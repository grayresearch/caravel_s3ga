VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO s3ga_proj
  CLASS BLOCK ;
  FOREIGN s3ga_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 1196.000 28.430 1200.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 1196.000 332.030 1200.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 1196.000 362.390 1200.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 1196.000 392.750 1200.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 1196.000 423.110 1200.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 1196.000 453.470 1200.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 1196.000 483.830 1200.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 1196.000 514.190 1200.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 1196.000 544.550 1200.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 1196.000 574.910 1200.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 1196.000 605.270 1200.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 1196.000 58.790 1200.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 1196.000 635.630 1200.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 1196.000 665.990 1200.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 1196.000 696.350 1200.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 1196.000 726.710 1200.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 1196.000 757.070 1200.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 1196.000 787.430 1200.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 1196.000 817.790 1200.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.870 1196.000 848.150 1200.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.230 1196.000 878.510 1200.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 1196.000 908.870 1200.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 1196.000 89.150 1200.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.950 1196.000 939.230 1200.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 1196.000 969.590 1200.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 1196.000 999.950 1200.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.030 1196.000 1030.310 1200.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.390 1196.000 1060.670 1200.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.750 1196.000 1091.030 1200.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 1196.000 1121.390 1200.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.470 1196.000 1151.750 1200.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1196.000 119.510 1200.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 1196.000 149.870 1200.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 1196.000 180.230 1200.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 1196.000 210.590 1200.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 1196.000 240.950 1200.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 1196.000 271.310 1200.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 1196.000 301.670 1200.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 1196.000 38.550 1200.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 1196.000 342.150 1200.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 1196.000 372.510 1200.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 1196.000 402.870 1200.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 1196.000 433.230 1200.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 1196.000 463.590 1200.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 1196.000 493.950 1200.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 1196.000 524.310 1200.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 1196.000 554.670 1200.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 1196.000 585.030 1200.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 1196.000 615.390 1200.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 1196.000 68.910 1200.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 1196.000 645.750 1200.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 1196.000 676.110 1200.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 1196.000 706.470 1200.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 1196.000 736.830 1200.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 1196.000 767.190 1200.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 1196.000 797.550 1200.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 1196.000 827.910 1200.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 1196.000 858.270 1200.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 1196.000 888.630 1200.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.710 1196.000 918.990 1200.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 1196.000 99.270 1200.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 1196.000 949.350 1200.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 1196.000 979.710 1200.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 1196.000 1010.070 1200.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 1196.000 1040.430 1200.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.510 1196.000 1070.790 1200.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.870 1196.000 1101.150 1200.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.230 1196.000 1131.510 1200.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.590 1196.000 1161.870 1200.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 1196.000 129.630 1200.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 1196.000 159.990 1200.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 1196.000 190.350 1200.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 1196.000 220.710 1200.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 1196.000 251.070 1200.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 1196.000 281.430 1200.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 1196.000 311.790 1200.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1196.000 48.670 1200.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 1196.000 352.270 1200.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 1196.000 382.630 1200.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 1196.000 412.990 1200.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 1196.000 443.350 1200.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 1196.000 473.710 1200.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 1196.000 504.070 1200.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 1196.000 534.430 1200.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 1196.000 564.790 1200.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 1196.000 595.150 1200.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 1196.000 625.510 1200.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 1196.000 79.030 1200.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 1196.000 655.870 1200.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 1196.000 686.230 1200.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 1196.000 716.590 1200.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 1196.000 746.950 1200.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 1196.000 777.310 1200.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 1196.000 807.670 1200.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 1196.000 838.030 1200.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 1196.000 868.390 1200.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 1196.000 898.750 1200.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 1196.000 929.110 1200.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 1196.000 109.390 1200.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 1196.000 959.470 1200.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 1196.000 989.830 1200.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.910 1196.000 1020.190 1200.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 1196.000 1050.550 1200.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 1196.000 1080.910 1200.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 1196.000 1111.270 1200.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 1196.000 1141.630 1200.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.710 1196.000 1171.990 1200.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 1196.000 139.750 1200.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 1196.000 170.110 1200.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 1196.000 200.470 1200.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 1196.000 230.830 1200.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 1196.000 261.190 1200.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 1196.000 291.550 1200.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 1196.000 321.910 1200.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 0.000 966.830 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.450 0.000 973.730 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 0.000 994.430 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.050 0.000 1001.330 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.850 0.000 1015.130 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.750 0.000 1022.030 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 0.000 1028.930 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.550 0.000 1035.830 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.450 0.000 1042.730 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.350 0.000 1049.630 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.150 0.000 1063.430 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 0.000 1070.330 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 0.000 1077.230 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.850 0.000 1084.130 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.750 0.000 1091.030 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.650 0.000 1097.930 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.450 0.000 1111.730 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.350 0.000 1118.630 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.250 0.000 1125.530 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.150 0.000 1132.430 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.050 0.000 1139.330 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 0.000 1146.230 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 0.000 635.630 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 0.000 642.530 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.950 0.000 663.230 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 0.000 746.030 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 0.000 759.830 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 0.000 801.230 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.650 0.000 821.930 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 0.000 835.730 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 0.000 842.630 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.250 0.000 849.530 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 0.000 856.430 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 0.000 870.230 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850 0.000 877.130 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.750 0.000 884.030 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.650 0.000 890.930 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.450 0.000 904.730 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 0.000 918.530 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.150 0.000 925.430 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.950 0.000 939.230 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.850 0.000 946.130 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 0.000 953.030 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 0.000 969.130 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 0.000 989.830 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 0.000 996.730 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.350 0.000 1003.630 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 0.000 1010.530 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 0.000 1017.430 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 0.000 1031.230 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 0.000 1038.130 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 0.000 1045.030 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 0.000 1051.930 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 0.000 1058.830 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 0.000 1065.730 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 0.000 1079.530 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 0.000 1086.430 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 0.000 1093.330 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.950 0.000 1100.230 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 0.000 1107.130 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.750 0.000 1114.030 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.550 0.000 1127.830 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 0.000 1141.630 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.250 0.000 1148.530 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.150 0.000 1155.430 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 0.000 651.730 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 0.000 658.630 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 0.000 672.430 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 0.000 755.230 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 0.000 762.130 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 0.000 796.630 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 0.000 803.530 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 0.000 824.230 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 0.000 838.030 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 0.000 844.930 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.550 0.000 851.830 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 0.000 858.730 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 0.000 865.630 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 0.000 886.330 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 0.000 893.230 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 0.000 900.130 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 0.000 907.030 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 0.000 920.830 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 0.000 934.630 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 0.000 941.530 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 0.000 948.430 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.950 0.000 962.230 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.150 0.000 971.430 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.050 0.000 978.330 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.650 0.000 1005.930 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 0.000 1012.830 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.450 0.000 1019.730 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 0.000 1026.630 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 0.000 1033.530 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 0.000 1047.330 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 0.000 1054.230 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.850 0.000 1061.130 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.750 0.000 1068.030 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.650 0.000 1074.930 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.550 0.000 1081.830 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 0.000 1095.630 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 0.000 1102.530 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 0.000 1109.430 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.050 0.000 1116.330 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.950 0.000 1123.230 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.850 0.000 1130.130 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.650 0.000 1143.930 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.550 0.000 1150.830 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 0.000 1157.730 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 0.000 598.830 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 0.000 681.630 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 0.000 695.430 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 0.000 736.830 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 0.000 743.730 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 0.000 764.430 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 0.000 771.330 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 0.000 792.030 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.350 0.000 819.630 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 0.000 833.430 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 0.000 840.330 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 0.000 854.130 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 0.000 874.830 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.150 0.000 902.430 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050 0.000 909.330 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 0.000 916.230 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.850 0.000 923.130 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 0.000 930.030 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.450 0.000 950.730 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 0.000 957.630 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.250 0.000 964.530 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.750 0.000 1160.030 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.050 0.000 1162.330 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.650 0.000 1166.930 4.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1188.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1188.880 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 5.330 1187.225 1194.350 1188.830 ;
        RECT 5.330 1181.785 1194.350 1184.615 ;
        RECT 5.330 1176.345 1194.350 1179.175 ;
        RECT 5.330 1170.905 1194.350 1173.735 ;
        RECT 5.330 1165.465 1194.350 1168.295 ;
        RECT 5.330 1160.025 1194.350 1162.855 ;
        RECT 5.330 1154.585 1194.350 1157.415 ;
        RECT 5.330 1149.145 1194.350 1151.975 ;
        RECT 5.330 1143.705 1194.350 1146.535 ;
        RECT 5.330 1138.265 1194.350 1141.095 ;
        RECT 5.330 1132.825 1194.350 1135.655 ;
        RECT 5.330 1127.385 1194.350 1130.215 ;
        RECT 5.330 1121.945 1194.350 1124.775 ;
        RECT 5.330 1116.505 1194.350 1119.335 ;
        RECT 5.330 1111.065 1194.350 1113.895 ;
        RECT 5.330 1105.625 1194.350 1108.455 ;
        RECT 5.330 1100.185 1194.350 1103.015 ;
        RECT 5.330 1094.745 1194.350 1097.575 ;
        RECT 5.330 1089.305 1194.350 1092.135 ;
        RECT 5.330 1083.865 1194.350 1086.695 ;
        RECT 5.330 1078.425 1194.350 1081.255 ;
        RECT 5.330 1072.985 1194.350 1075.815 ;
        RECT 5.330 1067.545 1194.350 1070.375 ;
        RECT 5.330 1062.105 1194.350 1064.935 ;
        RECT 5.330 1056.665 1194.350 1059.495 ;
        RECT 5.330 1051.225 1194.350 1054.055 ;
        RECT 5.330 1045.785 1194.350 1048.615 ;
        RECT 5.330 1040.345 1194.350 1043.175 ;
        RECT 5.330 1034.905 1194.350 1037.735 ;
        RECT 5.330 1029.465 1194.350 1032.295 ;
        RECT 5.330 1024.025 1194.350 1026.855 ;
        RECT 5.330 1018.585 1194.350 1021.415 ;
        RECT 5.330 1013.145 1194.350 1015.975 ;
        RECT 5.330 1007.705 1194.350 1010.535 ;
        RECT 5.330 1002.265 1194.350 1005.095 ;
        RECT 5.330 996.825 1194.350 999.655 ;
        RECT 5.330 991.385 1194.350 994.215 ;
        RECT 5.330 985.945 1194.350 988.775 ;
        RECT 5.330 980.505 1194.350 983.335 ;
        RECT 5.330 975.065 1194.350 977.895 ;
        RECT 5.330 969.625 1194.350 972.455 ;
        RECT 5.330 964.185 1194.350 967.015 ;
        RECT 5.330 958.745 1194.350 961.575 ;
        RECT 5.330 953.305 1194.350 956.135 ;
        RECT 5.330 947.865 1194.350 950.695 ;
        RECT 5.330 942.425 1194.350 945.255 ;
        RECT 5.330 936.985 1194.350 939.815 ;
        RECT 5.330 931.545 1194.350 934.375 ;
        RECT 5.330 926.105 1194.350 928.935 ;
        RECT 5.330 920.665 1194.350 923.495 ;
        RECT 5.330 915.225 1194.350 918.055 ;
        RECT 5.330 909.785 1194.350 912.615 ;
        RECT 5.330 904.345 1194.350 907.175 ;
        RECT 5.330 898.905 1194.350 901.735 ;
        RECT 5.330 893.465 1194.350 896.295 ;
        RECT 5.330 888.025 1194.350 890.855 ;
        RECT 5.330 882.585 1194.350 885.415 ;
        RECT 5.330 877.145 1194.350 879.975 ;
        RECT 5.330 871.705 1194.350 874.535 ;
        RECT 5.330 866.265 1194.350 869.095 ;
        RECT 5.330 860.825 1194.350 863.655 ;
        RECT 5.330 855.385 1194.350 858.215 ;
        RECT 5.330 849.945 1194.350 852.775 ;
        RECT 5.330 844.505 1194.350 847.335 ;
        RECT 5.330 839.065 1194.350 841.895 ;
        RECT 5.330 833.625 1194.350 836.455 ;
        RECT 5.330 828.185 1194.350 831.015 ;
        RECT 5.330 822.745 1194.350 825.575 ;
        RECT 5.330 817.305 1194.350 820.135 ;
        RECT 5.330 811.865 1194.350 814.695 ;
        RECT 5.330 806.425 1194.350 809.255 ;
        RECT 5.330 800.985 1194.350 803.815 ;
        RECT 5.330 795.545 1194.350 798.375 ;
        RECT 5.330 790.105 1194.350 792.935 ;
        RECT 5.330 784.665 1194.350 787.495 ;
        RECT 5.330 779.225 1194.350 782.055 ;
        RECT 5.330 773.785 1194.350 776.615 ;
        RECT 5.330 768.345 1194.350 771.175 ;
        RECT 5.330 762.905 1194.350 765.735 ;
        RECT 5.330 757.465 1194.350 760.295 ;
        RECT 5.330 752.025 1194.350 754.855 ;
        RECT 5.330 746.585 1194.350 749.415 ;
        RECT 5.330 741.145 1194.350 743.975 ;
        RECT 5.330 735.705 1194.350 738.535 ;
        RECT 5.330 730.265 1194.350 733.095 ;
        RECT 5.330 724.825 1194.350 727.655 ;
        RECT 5.330 719.385 1194.350 722.215 ;
        RECT 5.330 713.945 1194.350 716.775 ;
        RECT 5.330 708.505 1194.350 711.335 ;
        RECT 5.330 703.065 1194.350 705.895 ;
        RECT 5.330 697.625 1194.350 700.455 ;
        RECT 5.330 692.185 1194.350 695.015 ;
        RECT 5.330 686.745 1194.350 689.575 ;
        RECT 5.330 681.305 1194.350 684.135 ;
        RECT 5.330 675.865 1194.350 678.695 ;
        RECT 5.330 670.425 1194.350 673.255 ;
        RECT 5.330 664.985 1194.350 667.815 ;
        RECT 5.330 659.545 1194.350 662.375 ;
        RECT 5.330 654.105 1194.350 656.935 ;
        RECT 5.330 648.665 1194.350 651.495 ;
        RECT 5.330 643.225 1194.350 646.055 ;
        RECT 5.330 637.785 1194.350 640.615 ;
        RECT 5.330 632.345 1194.350 635.175 ;
        RECT 5.330 626.905 1194.350 629.735 ;
        RECT 5.330 621.465 1194.350 624.295 ;
        RECT 5.330 616.025 1194.350 618.855 ;
        RECT 5.330 610.585 1194.350 613.415 ;
        RECT 5.330 605.145 1194.350 607.975 ;
        RECT 5.330 599.705 1194.350 602.535 ;
        RECT 5.330 594.265 1194.350 597.095 ;
        RECT 5.330 588.825 1194.350 591.655 ;
        RECT 5.330 583.385 1194.350 586.215 ;
        RECT 5.330 577.945 1194.350 580.775 ;
        RECT 5.330 572.505 1194.350 575.335 ;
        RECT 5.330 567.065 1194.350 569.895 ;
        RECT 5.330 561.625 1194.350 564.455 ;
        RECT 5.330 556.185 1194.350 559.015 ;
        RECT 5.330 550.745 1194.350 553.575 ;
        RECT 5.330 545.305 1194.350 548.135 ;
        RECT 5.330 539.865 1194.350 542.695 ;
        RECT 5.330 534.425 1194.350 537.255 ;
        RECT 5.330 528.985 1194.350 531.815 ;
        RECT 5.330 523.545 1194.350 526.375 ;
        RECT 5.330 518.105 1194.350 520.935 ;
        RECT 5.330 512.665 1194.350 515.495 ;
        RECT 5.330 507.225 1194.350 510.055 ;
        RECT 5.330 501.785 1194.350 504.615 ;
        RECT 5.330 496.345 1194.350 499.175 ;
        RECT 5.330 490.905 1194.350 493.735 ;
        RECT 5.330 485.465 1194.350 488.295 ;
        RECT 5.330 480.025 1194.350 482.855 ;
        RECT 5.330 474.585 1194.350 477.415 ;
        RECT 5.330 469.145 1194.350 471.975 ;
        RECT 5.330 463.705 1194.350 466.535 ;
        RECT 5.330 458.265 1194.350 461.095 ;
        RECT 5.330 452.825 1194.350 455.655 ;
        RECT 5.330 447.385 1194.350 450.215 ;
        RECT 5.330 441.945 1194.350 444.775 ;
        RECT 5.330 436.505 1194.350 439.335 ;
        RECT 5.330 431.065 1194.350 433.895 ;
        RECT 5.330 425.625 1194.350 428.455 ;
        RECT 5.330 420.185 1194.350 423.015 ;
        RECT 5.330 414.745 1194.350 417.575 ;
        RECT 5.330 409.305 1194.350 412.135 ;
        RECT 5.330 403.865 1194.350 406.695 ;
        RECT 5.330 398.425 1194.350 401.255 ;
        RECT 5.330 392.985 1194.350 395.815 ;
        RECT 5.330 387.545 1194.350 390.375 ;
        RECT 5.330 382.105 1194.350 384.935 ;
        RECT 5.330 376.665 1194.350 379.495 ;
        RECT 5.330 371.225 1194.350 374.055 ;
        RECT 5.330 365.785 1194.350 368.615 ;
        RECT 5.330 360.345 1194.350 363.175 ;
        RECT 5.330 354.905 1194.350 357.735 ;
        RECT 5.330 349.465 1194.350 352.295 ;
        RECT 5.330 344.025 1194.350 346.855 ;
        RECT 5.330 338.585 1194.350 341.415 ;
        RECT 5.330 333.145 1194.350 335.975 ;
        RECT 5.330 327.705 1194.350 330.535 ;
        RECT 5.330 322.265 1194.350 325.095 ;
        RECT 5.330 316.825 1194.350 319.655 ;
        RECT 5.330 311.385 1194.350 314.215 ;
        RECT 5.330 305.945 1194.350 308.775 ;
        RECT 5.330 300.505 1194.350 303.335 ;
        RECT 5.330 295.065 1194.350 297.895 ;
        RECT 5.330 289.625 1194.350 292.455 ;
        RECT 5.330 284.185 1194.350 287.015 ;
        RECT 5.330 278.745 1194.350 281.575 ;
        RECT 5.330 273.305 1194.350 276.135 ;
        RECT 5.330 267.865 1194.350 270.695 ;
        RECT 5.330 262.425 1194.350 265.255 ;
        RECT 5.330 256.985 1194.350 259.815 ;
        RECT 5.330 251.545 1194.350 254.375 ;
        RECT 5.330 246.105 1194.350 248.935 ;
        RECT 5.330 240.665 1194.350 243.495 ;
        RECT 5.330 235.225 1194.350 238.055 ;
        RECT 5.330 229.785 1194.350 232.615 ;
        RECT 5.330 224.345 1194.350 227.175 ;
        RECT 5.330 218.905 1194.350 221.735 ;
        RECT 5.330 213.465 1194.350 216.295 ;
        RECT 5.330 208.025 1194.350 210.855 ;
        RECT 5.330 202.585 1194.350 205.415 ;
        RECT 5.330 197.145 1194.350 199.975 ;
        RECT 5.330 191.705 1194.350 194.535 ;
        RECT 5.330 186.265 1194.350 189.095 ;
        RECT 5.330 180.825 1194.350 183.655 ;
        RECT 5.330 175.385 1194.350 178.215 ;
        RECT 5.330 169.945 1194.350 172.775 ;
        RECT 5.330 164.505 1194.350 167.335 ;
        RECT 5.330 159.065 1194.350 161.895 ;
        RECT 5.330 153.625 1194.350 156.455 ;
        RECT 5.330 148.185 1194.350 151.015 ;
        RECT 5.330 142.745 1194.350 145.575 ;
        RECT 5.330 137.305 1194.350 140.135 ;
        RECT 5.330 131.865 1194.350 134.695 ;
        RECT 5.330 126.425 1194.350 129.255 ;
        RECT 5.330 120.985 1194.350 123.815 ;
        RECT 5.330 115.545 1194.350 118.375 ;
        RECT 5.330 110.105 1194.350 112.935 ;
        RECT 5.330 104.665 1194.350 107.495 ;
        RECT 5.330 99.225 1194.350 102.055 ;
        RECT 5.330 93.785 1194.350 96.615 ;
        RECT 5.330 88.345 1194.350 91.175 ;
        RECT 5.330 82.905 1194.350 85.735 ;
        RECT 5.330 77.465 1194.350 80.295 ;
        RECT 5.330 72.025 1194.350 74.855 ;
        RECT 5.330 66.585 1194.350 69.415 ;
        RECT 5.330 61.145 1194.350 63.975 ;
        RECT 5.330 55.705 1194.350 58.535 ;
        RECT 5.330 50.265 1194.350 53.095 ;
        RECT 5.330 44.825 1194.350 47.655 ;
        RECT 5.330 39.385 1194.350 42.215 ;
        RECT 5.330 33.945 1194.350 36.775 ;
        RECT 5.330 28.505 1194.350 31.335 ;
        RECT 5.330 23.065 1194.350 25.895 ;
        RECT 5.330 17.625 1194.350 20.455 ;
        RECT 5.330 12.185 1194.350 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 1188.725 ;
      LAYER met1 ;
        RECT 5.520 2.420 1194.160 1189.960 ;
      LAYER met2 ;
        RECT 7.920 1195.720 27.870 1196.530 ;
        RECT 28.710 1195.720 37.990 1196.530 ;
        RECT 38.830 1195.720 48.110 1196.530 ;
        RECT 48.950 1195.720 58.230 1196.530 ;
        RECT 59.070 1195.720 68.350 1196.530 ;
        RECT 69.190 1195.720 78.470 1196.530 ;
        RECT 79.310 1195.720 88.590 1196.530 ;
        RECT 89.430 1195.720 98.710 1196.530 ;
        RECT 99.550 1195.720 108.830 1196.530 ;
        RECT 109.670 1195.720 118.950 1196.530 ;
        RECT 119.790 1195.720 129.070 1196.530 ;
        RECT 129.910 1195.720 139.190 1196.530 ;
        RECT 140.030 1195.720 149.310 1196.530 ;
        RECT 150.150 1195.720 159.430 1196.530 ;
        RECT 160.270 1195.720 169.550 1196.530 ;
        RECT 170.390 1195.720 179.670 1196.530 ;
        RECT 180.510 1195.720 189.790 1196.530 ;
        RECT 190.630 1195.720 199.910 1196.530 ;
        RECT 200.750 1195.720 210.030 1196.530 ;
        RECT 210.870 1195.720 220.150 1196.530 ;
        RECT 220.990 1195.720 230.270 1196.530 ;
        RECT 231.110 1195.720 240.390 1196.530 ;
        RECT 241.230 1195.720 250.510 1196.530 ;
        RECT 251.350 1195.720 260.630 1196.530 ;
        RECT 261.470 1195.720 270.750 1196.530 ;
        RECT 271.590 1195.720 280.870 1196.530 ;
        RECT 281.710 1195.720 290.990 1196.530 ;
        RECT 291.830 1195.720 301.110 1196.530 ;
        RECT 301.950 1195.720 311.230 1196.530 ;
        RECT 312.070 1195.720 321.350 1196.530 ;
        RECT 322.190 1195.720 331.470 1196.530 ;
        RECT 332.310 1195.720 341.590 1196.530 ;
        RECT 342.430 1195.720 351.710 1196.530 ;
        RECT 352.550 1195.720 361.830 1196.530 ;
        RECT 362.670 1195.720 371.950 1196.530 ;
        RECT 372.790 1195.720 382.070 1196.530 ;
        RECT 382.910 1195.720 392.190 1196.530 ;
        RECT 393.030 1195.720 402.310 1196.530 ;
        RECT 403.150 1195.720 412.430 1196.530 ;
        RECT 413.270 1195.720 422.550 1196.530 ;
        RECT 423.390 1195.720 432.670 1196.530 ;
        RECT 433.510 1195.720 442.790 1196.530 ;
        RECT 443.630 1195.720 452.910 1196.530 ;
        RECT 453.750 1195.720 463.030 1196.530 ;
        RECT 463.870 1195.720 473.150 1196.530 ;
        RECT 473.990 1195.720 483.270 1196.530 ;
        RECT 484.110 1195.720 493.390 1196.530 ;
        RECT 494.230 1195.720 503.510 1196.530 ;
        RECT 504.350 1195.720 513.630 1196.530 ;
        RECT 514.470 1195.720 523.750 1196.530 ;
        RECT 524.590 1195.720 533.870 1196.530 ;
        RECT 534.710 1195.720 543.990 1196.530 ;
        RECT 544.830 1195.720 554.110 1196.530 ;
        RECT 554.950 1195.720 564.230 1196.530 ;
        RECT 565.070 1195.720 574.350 1196.530 ;
        RECT 575.190 1195.720 584.470 1196.530 ;
        RECT 585.310 1195.720 594.590 1196.530 ;
        RECT 595.430 1195.720 604.710 1196.530 ;
        RECT 605.550 1195.720 614.830 1196.530 ;
        RECT 615.670 1195.720 624.950 1196.530 ;
        RECT 625.790 1195.720 635.070 1196.530 ;
        RECT 635.910 1195.720 645.190 1196.530 ;
        RECT 646.030 1195.720 655.310 1196.530 ;
        RECT 656.150 1195.720 665.430 1196.530 ;
        RECT 666.270 1195.720 675.550 1196.530 ;
        RECT 676.390 1195.720 685.670 1196.530 ;
        RECT 686.510 1195.720 695.790 1196.530 ;
        RECT 696.630 1195.720 705.910 1196.530 ;
        RECT 706.750 1195.720 716.030 1196.530 ;
        RECT 716.870 1195.720 726.150 1196.530 ;
        RECT 726.990 1195.720 736.270 1196.530 ;
        RECT 737.110 1195.720 746.390 1196.530 ;
        RECT 747.230 1195.720 756.510 1196.530 ;
        RECT 757.350 1195.720 766.630 1196.530 ;
        RECT 767.470 1195.720 776.750 1196.530 ;
        RECT 777.590 1195.720 786.870 1196.530 ;
        RECT 787.710 1195.720 796.990 1196.530 ;
        RECT 797.830 1195.720 807.110 1196.530 ;
        RECT 807.950 1195.720 817.230 1196.530 ;
        RECT 818.070 1195.720 827.350 1196.530 ;
        RECT 828.190 1195.720 837.470 1196.530 ;
        RECT 838.310 1195.720 847.590 1196.530 ;
        RECT 848.430 1195.720 857.710 1196.530 ;
        RECT 858.550 1195.720 867.830 1196.530 ;
        RECT 868.670 1195.720 877.950 1196.530 ;
        RECT 878.790 1195.720 888.070 1196.530 ;
        RECT 888.910 1195.720 898.190 1196.530 ;
        RECT 899.030 1195.720 908.310 1196.530 ;
        RECT 909.150 1195.720 918.430 1196.530 ;
        RECT 919.270 1195.720 928.550 1196.530 ;
        RECT 929.390 1195.720 938.670 1196.530 ;
        RECT 939.510 1195.720 948.790 1196.530 ;
        RECT 949.630 1195.720 958.910 1196.530 ;
        RECT 959.750 1195.720 969.030 1196.530 ;
        RECT 969.870 1195.720 979.150 1196.530 ;
        RECT 979.990 1195.720 989.270 1196.530 ;
        RECT 990.110 1195.720 999.390 1196.530 ;
        RECT 1000.230 1195.720 1009.510 1196.530 ;
        RECT 1010.350 1195.720 1019.630 1196.530 ;
        RECT 1020.470 1195.720 1029.750 1196.530 ;
        RECT 1030.590 1195.720 1039.870 1196.530 ;
        RECT 1040.710 1195.720 1049.990 1196.530 ;
        RECT 1050.830 1195.720 1060.110 1196.530 ;
        RECT 1060.950 1195.720 1070.230 1196.530 ;
        RECT 1071.070 1195.720 1080.350 1196.530 ;
        RECT 1081.190 1195.720 1090.470 1196.530 ;
        RECT 1091.310 1195.720 1100.590 1196.530 ;
        RECT 1101.430 1195.720 1110.710 1196.530 ;
        RECT 1111.550 1195.720 1120.830 1196.530 ;
        RECT 1121.670 1195.720 1130.950 1196.530 ;
        RECT 1131.790 1195.720 1141.070 1196.530 ;
        RECT 1141.910 1195.720 1151.190 1196.530 ;
        RECT 1152.030 1195.720 1161.310 1196.530 ;
        RECT 1162.150 1195.720 1171.430 1196.530 ;
        RECT 1172.270 1195.720 1192.220 1196.530 ;
        RECT 7.920 4.280 1192.220 1195.720 ;
        RECT 7.920 2.390 32.470 4.280 ;
        RECT 33.310 2.390 34.770 4.280 ;
        RECT 35.610 2.390 37.070 4.280 ;
        RECT 37.910 2.390 39.370 4.280 ;
        RECT 40.210 2.390 41.670 4.280 ;
        RECT 42.510 2.390 43.970 4.280 ;
        RECT 44.810 2.390 46.270 4.280 ;
        RECT 47.110 2.390 48.570 4.280 ;
        RECT 49.410 2.390 50.870 4.280 ;
        RECT 51.710 2.390 53.170 4.280 ;
        RECT 54.010 2.390 55.470 4.280 ;
        RECT 56.310 2.390 57.770 4.280 ;
        RECT 58.610 2.390 60.070 4.280 ;
        RECT 60.910 2.390 62.370 4.280 ;
        RECT 63.210 2.390 64.670 4.280 ;
        RECT 65.510 2.390 66.970 4.280 ;
        RECT 67.810 2.390 69.270 4.280 ;
        RECT 70.110 2.390 71.570 4.280 ;
        RECT 72.410 2.390 73.870 4.280 ;
        RECT 74.710 2.390 76.170 4.280 ;
        RECT 77.010 2.390 78.470 4.280 ;
        RECT 79.310 2.390 80.770 4.280 ;
        RECT 81.610 2.390 83.070 4.280 ;
        RECT 83.910 2.390 85.370 4.280 ;
        RECT 86.210 2.390 87.670 4.280 ;
        RECT 88.510 2.390 89.970 4.280 ;
        RECT 90.810 2.390 92.270 4.280 ;
        RECT 93.110 2.390 94.570 4.280 ;
        RECT 95.410 2.390 96.870 4.280 ;
        RECT 97.710 2.390 99.170 4.280 ;
        RECT 100.010 2.390 101.470 4.280 ;
        RECT 102.310 2.390 103.770 4.280 ;
        RECT 104.610 2.390 106.070 4.280 ;
        RECT 106.910 2.390 108.370 4.280 ;
        RECT 109.210 2.390 110.670 4.280 ;
        RECT 111.510 2.390 112.970 4.280 ;
        RECT 113.810 2.390 115.270 4.280 ;
        RECT 116.110 2.390 117.570 4.280 ;
        RECT 118.410 2.390 119.870 4.280 ;
        RECT 120.710 2.390 122.170 4.280 ;
        RECT 123.010 2.390 124.470 4.280 ;
        RECT 125.310 2.390 126.770 4.280 ;
        RECT 127.610 2.390 129.070 4.280 ;
        RECT 129.910 2.390 131.370 4.280 ;
        RECT 132.210 2.390 133.670 4.280 ;
        RECT 134.510 2.390 135.970 4.280 ;
        RECT 136.810 2.390 138.270 4.280 ;
        RECT 139.110 2.390 140.570 4.280 ;
        RECT 141.410 2.390 142.870 4.280 ;
        RECT 143.710 2.390 145.170 4.280 ;
        RECT 146.010 2.390 147.470 4.280 ;
        RECT 148.310 2.390 149.770 4.280 ;
        RECT 150.610 2.390 152.070 4.280 ;
        RECT 152.910 2.390 154.370 4.280 ;
        RECT 155.210 2.390 156.670 4.280 ;
        RECT 157.510 2.390 158.970 4.280 ;
        RECT 159.810 2.390 161.270 4.280 ;
        RECT 162.110 2.390 163.570 4.280 ;
        RECT 164.410 2.390 165.870 4.280 ;
        RECT 166.710 2.390 168.170 4.280 ;
        RECT 169.010 2.390 170.470 4.280 ;
        RECT 171.310 2.390 172.770 4.280 ;
        RECT 173.610 2.390 175.070 4.280 ;
        RECT 175.910 2.390 177.370 4.280 ;
        RECT 178.210 2.390 179.670 4.280 ;
        RECT 180.510 2.390 181.970 4.280 ;
        RECT 182.810 2.390 184.270 4.280 ;
        RECT 185.110 2.390 186.570 4.280 ;
        RECT 187.410 2.390 188.870 4.280 ;
        RECT 189.710 2.390 191.170 4.280 ;
        RECT 192.010 2.390 193.470 4.280 ;
        RECT 194.310 2.390 195.770 4.280 ;
        RECT 196.610 2.390 198.070 4.280 ;
        RECT 198.910 2.390 200.370 4.280 ;
        RECT 201.210 2.390 202.670 4.280 ;
        RECT 203.510 2.390 204.970 4.280 ;
        RECT 205.810 2.390 207.270 4.280 ;
        RECT 208.110 2.390 209.570 4.280 ;
        RECT 210.410 2.390 211.870 4.280 ;
        RECT 212.710 2.390 214.170 4.280 ;
        RECT 215.010 2.390 216.470 4.280 ;
        RECT 217.310 2.390 218.770 4.280 ;
        RECT 219.610 2.390 221.070 4.280 ;
        RECT 221.910 2.390 223.370 4.280 ;
        RECT 224.210 2.390 225.670 4.280 ;
        RECT 226.510 2.390 227.970 4.280 ;
        RECT 228.810 2.390 230.270 4.280 ;
        RECT 231.110 2.390 232.570 4.280 ;
        RECT 233.410 2.390 234.870 4.280 ;
        RECT 235.710 2.390 237.170 4.280 ;
        RECT 238.010 2.390 239.470 4.280 ;
        RECT 240.310 2.390 241.770 4.280 ;
        RECT 242.610 2.390 244.070 4.280 ;
        RECT 244.910 2.390 246.370 4.280 ;
        RECT 247.210 2.390 248.670 4.280 ;
        RECT 249.510 2.390 250.970 4.280 ;
        RECT 251.810 2.390 253.270 4.280 ;
        RECT 254.110 2.390 255.570 4.280 ;
        RECT 256.410 2.390 257.870 4.280 ;
        RECT 258.710 2.390 260.170 4.280 ;
        RECT 261.010 2.390 262.470 4.280 ;
        RECT 263.310 2.390 264.770 4.280 ;
        RECT 265.610 2.390 267.070 4.280 ;
        RECT 267.910 2.390 269.370 4.280 ;
        RECT 270.210 2.390 271.670 4.280 ;
        RECT 272.510 2.390 273.970 4.280 ;
        RECT 274.810 2.390 276.270 4.280 ;
        RECT 277.110 2.390 278.570 4.280 ;
        RECT 279.410 2.390 280.870 4.280 ;
        RECT 281.710 2.390 283.170 4.280 ;
        RECT 284.010 2.390 285.470 4.280 ;
        RECT 286.310 2.390 287.770 4.280 ;
        RECT 288.610 2.390 290.070 4.280 ;
        RECT 290.910 2.390 292.370 4.280 ;
        RECT 293.210 2.390 294.670 4.280 ;
        RECT 295.510 2.390 296.970 4.280 ;
        RECT 297.810 2.390 299.270 4.280 ;
        RECT 300.110 2.390 301.570 4.280 ;
        RECT 302.410 2.390 303.870 4.280 ;
        RECT 304.710 2.390 306.170 4.280 ;
        RECT 307.010 2.390 308.470 4.280 ;
        RECT 309.310 2.390 310.770 4.280 ;
        RECT 311.610 2.390 313.070 4.280 ;
        RECT 313.910 2.390 315.370 4.280 ;
        RECT 316.210 2.390 317.670 4.280 ;
        RECT 318.510 2.390 319.970 4.280 ;
        RECT 320.810 2.390 322.270 4.280 ;
        RECT 323.110 2.390 324.570 4.280 ;
        RECT 325.410 2.390 326.870 4.280 ;
        RECT 327.710 2.390 329.170 4.280 ;
        RECT 330.010 2.390 331.470 4.280 ;
        RECT 332.310 2.390 333.770 4.280 ;
        RECT 334.610 2.390 336.070 4.280 ;
        RECT 336.910 2.390 338.370 4.280 ;
        RECT 339.210 2.390 340.670 4.280 ;
        RECT 341.510 2.390 342.970 4.280 ;
        RECT 343.810 2.390 345.270 4.280 ;
        RECT 346.110 2.390 347.570 4.280 ;
        RECT 348.410 2.390 349.870 4.280 ;
        RECT 350.710 2.390 352.170 4.280 ;
        RECT 353.010 2.390 354.470 4.280 ;
        RECT 355.310 2.390 356.770 4.280 ;
        RECT 357.610 2.390 359.070 4.280 ;
        RECT 359.910 2.390 361.370 4.280 ;
        RECT 362.210 2.390 363.670 4.280 ;
        RECT 364.510 2.390 365.970 4.280 ;
        RECT 366.810 2.390 368.270 4.280 ;
        RECT 369.110 2.390 370.570 4.280 ;
        RECT 371.410 2.390 372.870 4.280 ;
        RECT 373.710 2.390 375.170 4.280 ;
        RECT 376.010 2.390 377.470 4.280 ;
        RECT 378.310 2.390 379.770 4.280 ;
        RECT 380.610 2.390 382.070 4.280 ;
        RECT 382.910 2.390 384.370 4.280 ;
        RECT 385.210 2.390 386.670 4.280 ;
        RECT 387.510 2.390 388.970 4.280 ;
        RECT 389.810 2.390 391.270 4.280 ;
        RECT 392.110 2.390 393.570 4.280 ;
        RECT 394.410 2.390 395.870 4.280 ;
        RECT 396.710 2.390 398.170 4.280 ;
        RECT 399.010 2.390 400.470 4.280 ;
        RECT 401.310 2.390 402.770 4.280 ;
        RECT 403.610 2.390 405.070 4.280 ;
        RECT 405.910 2.390 407.370 4.280 ;
        RECT 408.210 2.390 409.670 4.280 ;
        RECT 410.510 2.390 411.970 4.280 ;
        RECT 412.810 2.390 414.270 4.280 ;
        RECT 415.110 2.390 416.570 4.280 ;
        RECT 417.410 2.390 418.870 4.280 ;
        RECT 419.710 2.390 421.170 4.280 ;
        RECT 422.010 2.390 423.470 4.280 ;
        RECT 424.310 2.390 425.770 4.280 ;
        RECT 426.610 2.390 428.070 4.280 ;
        RECT 428.910 2.390 430.370 4.280 ;
        RECT 431.210 2.390 432.670 4.280 ;
        RECT 433.510 2.390 434.970 4.280 ;
        RECT 435.810 2.390 437.270 4.280 ;
        RECT 438.110 2.390 439.570 4.280 ;
        RECT 440.410 2.390 441.870 4.280 ;
        RECT 442.710 2.390 444.170 4.280 ;
        RECT 445.010 2.390 446.470 4.280 ;
        RECT 447.310 2.390 448.770 4.280 ;
        RECT 449.610 2.390 451.070 4.280 ;
        RECT 451.910 2.390 453.370 4.280 ;
        RECT 454.210 2.390 455.670 4.280 ;
        RECT 456.510 2.390 457.970 4.280 ;
        RECT 458.810 2.390 460.270 4.280 ;
        RECT 461.110 2.390 462.570 4.280 ;
        RECT 463.410 2.390 464.870 4.280 ;
        RECT 465.710 2.390 467.170 4.280 ;
        RECT 468.010 2.390 469.470 4.280 ;
        RECT 470.310 2.390 471.770 4.280 ;
        RECT 472.610 2.390 474.070 4.280 ;
        RECT 474.910 2.390 476.370 4.280 ;
        RECT 477.210 2.390 478.670 4.280 ;
        RECT 479.510 2.390 480.970 4.280 ;
        RECT 481.810 2.390 483.270 4.280 ;
        RECT 484.110 2.390 485.570 4.280 ;
        RECT 486.410 2.390 487.870 4.280 ;
        RECT 488.710 2.390 490.170 4.280 ;
        RECT 491.010 2.390 492.470 4.280 ;
        RECT 493.310 2.390 494.770 4.280 ;
        RECT 495.610 2.390 497.070 4.280 ;
        RECT 497.910 2.390 499.370 4.280 ;
        RECT 500.210 2.390 501.670 4.280 ;
        RECT 502.510 2.390 503.970 4.280 ;
        RECT 504.810 2.390 506.270 4.280 ;
        RECT 507.110 2.390 508.570 4.280 ;
        RECT 509.410 2.390 510.870 4.280 ;
        RECT 511.710 2.390 513.170 4.280 ;
        RECT 514.010 2.390 515.470 4.280 ;
        RECT 516.310 2.390 517.770 4.280 ;
        RECT 518.610 2.390 520.070 4.280 ;
        RECT 520.910 2.390 522.370 4.280 ;
        RECT 523.210 2.390 524.670 4.280 ;
        RECT 525.510 2.390 526.970 4.280 ;
        RECT 527.810 2.390 529.270 4.280 ;
        RECT 530.110 2.390 531.570 4.280 ;
        RECT 532.410 2.390 533.870 4.280 ;
        RECT 534.710 2.390 536.170 4.280 ;
        RECT 537.010 2.390 538.470 4.280 ;
        RECT 539.310 2.390 540.770 4.280 ;
        RECT 541.610 2.390 543.070 4.280 ;
        RECT 543.910 2.390 545.370 4.280 ;
        RECT 546.210 2.390 547.670 4.280 ;
        RECT 548.510 2.390 549.970 4.280 ;
        RECT 550.810 2.390 552.270 4.280 ;
        RECT 553.110 2.390 554.570 4.280 ;
        RECT 555.410 2.390 556.870 4.280 ;
        RECT 557.710 2.390 559.170 4.280 ;
        RECT 560.010 2.390 561.470 4.280 ;
        RECT 562.310 2.390 563.770 4.280 ;
        RECT 564.610 2.390 566.070 4.280 ;
        RECT 566.910 2.390 568.370 4.280 ;
        RECT 569.210 2.390 570.670 4.280 ;
        RECT 571.510 2.390 572.970 4.280 ;
        RECT 573.810 2.390 575.270 4.280 ;
        RECT 576.110 2.390 577.570 4.280 ;
        RECT 578.410 2.390 579.870 4.280 ;
        RECT 580.710 2.390 582.170 4.280 ;
        RECT 583.010 2.390 584.470 4.280 ;
        RECT 585.310 2.390 586.770 4.280 ;
        RECT 587.610 2.390 589.070 4.280 ;
        RECT 589.910 2.390 591.370 4.280 ;
        RECT 592.210 2.390 593.670 4.280 ;
        RECT 594.510 2.390 595.970 4.280 ;
        RECT 596.810 2.390 598.270 4.280 ;
        RECT 599.110 2.390 600.570 4.280 ;
        RECT 601.410 2.390 602.870 4.280 ;
        RECT 603.710 2.390 605.170 4.280 ;
        RECT 606.010 2.390 607.470 4.280 ;
        RECT 608.310 2.390 609.770 4.280 ;
        RECT 610.610 2.390 612.070 4.280 ;
        RECT 612.910 2.390 614.370 4.280 ;
        RECT 615.210 2.390 616.670 4.280 ;
        RECT 617.510 2.390 618.970 4.280 ;
        RECT 619.810 2.390 621.270 4.280 ;
        RECT 622.110 2.390 623.570 4.280 ;
        RECT 624.410 2.390 625.870 4.280 ;
        RECT 626.710 2.390 628.170 4.280 ;
        RECT 629.010 2.390 630.470 4.280 ;
        RECT 631.310 2.390 632.770 4.280 ;
        RECT 633.610 2.390 635.070 4.280 ;
        RECT 635.910 2.390 637.370 4.280 ;
        RECT 638.210 2.390 639.670 4.280 ;
        RECT 640.510 2.390 641.970 4.280 ;
        RECT 642.810 2.390 644.270 4.280 ;
        RECT 645.110 2.390 646.570 4.280 ;
        RECT 647.410 2.390 648.870 4.280 ;
        RECT 649.710 2.390 651.170 4.280 ;
        RECT 652.010 2.390 653.470 4.280 ;
        RECT 654.310 2.390 655.770 4.280 ;
        RECT 656.610 2.390 658.070 4.280 ;
        RECT 658.910 2.390 660.370 4.280 ;
        RECT 661.210 2.390 662.670 4.280 ;
        RECT 663.510 2.390 664.970 4.280 ;
        RECT 665.810 2.390 667.270 4.280 ;
        RECT 668.110 2.390 669.570 4.280 ;
        RECT 670.410 2.390 671.870 4.280 ;
        RECT 672.710 2.390 674.170 4.280 ;
        RECT 675.010 2.390 676.470 4.280 ;
        RECT 677.310 2.390 678.770 4.280 ;
        RECT 679.610 2.390 681.070 4.280 ;
        RECT 681.910 2.390 683.370 4.280 ;
        RECT 684.210 2.390 685.670 4.280 ;
        RECT 686.510 2.390 687.970 4.280 ;
        RECT 688.810 2.390 690.270 4.280 ;
        RECT 691.110 2.390 692.570 4.280 ;
        RECT 693.410 2.390 694.870 4.280 ;
        RECT 695.710 2.390 697.170 4.280 ;
        RECT 698.010 2.390 699.470 4.280 ;
        RECT 700.310 2.390 701.770 4.280 ;
        RECT 702.610 2.390 704.070 4.280 ;
        RECT 704.910 2.390 706.370 4.280 ;
        RECT 707.210 2.390 708.670 4.280 ;
        RECT 709.510 2.390 710.970 4.280 ;
        RECT 711.810 2.390 713.270 4.280 ;
        RECT 714.110 2.390 715.570 4.280 ;
        RECT 716.410 2.390 717.870 4.280 ;
        RECT 718.710 2.390 720.170 4.280 ;
        RECT 721.010 2.390 722.470 4.280 ;
        RECT 723.310 2.390 724.770 4.280 ;
        RECT 725.610 2.390 727.070 4.280 ;
        RECT 727.910 2.390 729.370 4.280 ;
        RECT 730.210 2.390 731.670 4.280 ;
        RECT 732.510 2.390 733.970 4.280 ;
        RECT 734.810 2.390 736.270 4.280 ;
        RECT 737.110 2.390 738.570 4.280 ;
        RECT 739.410 2.390 740.870 4.280 ;
        RECT 741.710 2.390 743.170 4.280 ;
        RECT 744.010 2.390 745.470 4.280 ;
        RECT 746.310 2.390 747.770 4.280 ;
        RECT 748.610 2.390 750.070 4.280 ;
        RECT 750.910 2.390 752.370 4.280 ;
        RECT 753.210 2.390 754.670 4.280 ;
        RECT 755.510 2.390 756.970 4.280 ;
        RECT 757.810 2.390 759.270 4.280 ;
        RECT 760.110 2.390 761.570 4.280 ;
        RECT 762.410 2.390 763.870 4.280 ;
        RECT 764.710 2.390 766.170 4.280 ;
        RECT 767.010 2.390 768.470 4.280 ;
        RECT 769.310 2.390 770.770 4.280 ;
        RECT 771.610 2.390 773.070 4.280 ;
        RECT 773.910 2.390 775.370 4.280 ;
        RECT 776.210 2.390 777.670 4.280 ;
        RECT 778.510 2.390 779.970 4.280 ;
        RECT 780.810 2.390 782.270 4.280 ;
        RECT 783.110 2.390 784.570 4.280 ;
        RECT 785.410 2.390 786.870 4.280 ;
        RECT 787.710 2.390 789.170 4.280 ;
        RECT 790.010 2.390 791.470 4.280 ;
        RECT 792.310 2.390 793.770 4.280 ;
        RECT 794.610 2.390 796.070 4.280 ;
        RECT 796.910 2.390 798.370 4.280 ;
        RECT 799.210 2.390 800.670 4.280 ;
        RECT 801.510 2.390 802.970 4.280 ;
        RECT 803.810 2.390 805.270 4.280 ;
        RECT 806.110 2.390 807.570 4.280 ;
        RECT 808.410 2.390 809.870 4.280 ;
        RECT 810.710 2.390 812.170 4.280 ;
        RECT 813.010 2.390 814.470 4.280 ;
        RECT 815.310 2.390 816.770 4.280 ;
        RECT 817.610 2.390 819.070 4.280 ;
        RECT 819.910 2.390 821.370 4.280 ;
        RECT 822.210 2.390 823.670 4.280 ;
        RECT 824.510 2.390 825.970 4.280 ;
        RECT 826.810 2.390 828.270 4.280 ;
        RECT 829.110 2.390 830.570 4.280 ;
        RECT 831.410 2.390 832.870 4.280 ;
        RECT 833.710 2.390 835.170 4.280 ;
        RECT 836.010 2.390 837.470 4.280 ;
        RECT 838.310 2.390 839.770 4.280 ;
        RECT 840.610 2.390 842.070 4.280 ;
        RECT 842.910 2.390 844.370 4.280 ;
        RECT 845.210 2.390 846.670 4.280 ;
        RECT 847.510 2.390 848.970 4.280 ;
        RECT 849.810 2.390 851.270 4.280 ;
        RECT 852.110 2.390 853.570 4.280 ;
        RECT 854.410 2.390 855.870 4.280 ;
        RECT 856.710 2.390 858.170 4.280 ;
        RECT 859.010 2.390 860.470 4.280 ;
        RECT 861.310 2.390 862.770 4.280 ;
        RECT 863.610 2.390 865.070 4.280 ;
        RECT 865.910 2.390 867.370 4.280 ;
        RECT 868.210 2.390 869.670 4.280 ;
        RECT 870.510 2.390 871.970 4.280 ;
        RECT 872.810 2.390 874.270 4.280 ;
        RECT 875.110 2.390 876.570 4.280 ;
        RECT 877.410 2.390 878.870 4.280 ;
        RECT 879.710 2.390 881.170 4.280 ;
        RECT 882.010 2.390 883.470 4.280 ;
        RECT 884.310 2.390 885.770 4.280 ;
        RECT 886.610 2.390 888.070 4.280 ;
        RECT 888.910 2.390 890.370 4.280 ;
        RECT 891.210 2.390 892.670 4.280 ;
        RECT 893.510 2.390 894.970 4.280 ;
        RECT 895.810 2.390 897.270 4.280 ;
        RECT 898.110 2.390 899.570 4.280 ;
        RECT 900.410 2.390 901.870 4.280 ;
        RECT 902.710 2.390 904.170 4.280 ;
        RECT 905.010 2.390 906.470 4.280 ;
        RECT 907.310 2.390 908.770 4.280 ;
        RECT 909.610 2.390 911.070 4.280 ;
        RECT 911.910 2.390 913.370 4.280 ;
        RECT 914.210 2.390 915.670 4.280 ;
        RECT 916.510 2.390 917.970 4.280 ;
        RECT 918.810 2.390 920.270 4.280 ;
        RECT 921.110 2.390 922.570 4.280 ;
        RECT 923.410 2.390 924.870 4.280 ;
        RECT 925.710 2.390 927.170 4.280 ;
        RECT 928.010 2.390 929.470 4.280 ;
        RECT 930.310 2.390 931.770 4.280 ;
        RECT 932.610 2.390 934.070 4.280 ;
        RECT 934.910 2.390 936.370 4.280 ;
        RECT 937.210 2.390 938.670 4.280 ;
        RECT 939.510 2.390 940.970 4.280 ;
        RECT 941.810 2.390 943.270 4.280 ;
        RECT 944.110 2.390 945.570 4.280 ;
        RECT 946.410 2.390 947.870 4.280 ;
        RECT 948.710 2.390 950.170 4.280 ;
        RECT 951.010 2.390 952.470 4.280 ;
        RECT 953.310 2.390 954.770 4.280 ;
        RECT 955.610 2.390 957.070 4.280 ;
        RECT 957.910 2.390 959.370 4.280 ;
        RECT 960.210 2.390 961.670 4.280 ;
        RECT 962.510 2.390 963.970 4.280 ;
        RECT 964.810 2.390 966.270 4.280 ;
        RECT 967.110 2.390 968.570 4.280 ;
        RECT 969.410 2.390 970.870 4.280 ;
        RECT 971.710 2.390 973.170 4.280 ;
        RECT 974.010 2.390 975.470 4.280 ;
        RECT 976.310 2.390 977.770 4.280 ;
        RECT 978.610 2.390 980.070 4.280 ;
        RECT 980.910 2.390 982.370 4.280 ;
        RECT 983.210 2.390 984.670 4.280 ;
        RECT 985.510 2.390 986.970 4.280 ;
        RECT 987.810 2.390 989.270 4.280 ;
        RECT 990.110 2.390 991.570 4.280 ;
        RECT 992.410 2.390 993.870 4.280 ;
        RECT 994.710 2.390 996.170 4.280 ;
        RECT 997.010 2.390 998.470 4.280 ;
        RECT 999.310 2.390 1000.770 4.280 ;
        RECT 1001.610 2.390 1003.070 4.280 ;
        RECT 1003.910 2.390 1005.370 4.280 ;
        RECT 1006.210 2.390 1007.670 4.280 ;
        RECT 1008.510 2.390 1009.970 4.280 ;
        RECT 1010.810 2.390 1012.270 4.280 ;
        RECT 1013.110 2.390 1014.570 4.280 ;
        RECT 1015.410 2.390 1016.870 4.280 ;
        RECT 1017.710 2.390 1019.170 4.280 ;
        RECT 1020.010 2.390 1021.470 4.280 ;
        RECT 1022.310 2.390 1023.770 4.280 ;
        RECT 1024.610 2.390 1026.070 4.280 ;
        RECT 1026.910 2.390 1028.370 4.280 ;
        RECT 1029.210 2.390 1030.670 4.280 ;
        RECT 1031.510 2.390 1032.970 4.280 ;
        RECT 1033.810 2.390 1035.270 4.280 ;
        RECT 1036.110 2.390 1037.570 4.280 ;
        RECT 1038.410 2.390 1039.870 4.280 ;
        RECT 1040.710 2.390 1042.170 4.280 ;
        RECT 1043.010 2.390 1044.470 4.280 ;
        RECT 1045.310 2.390 1046.770 4.280 ;
        RECT 1047.610 2.390 1049.070 4.280 ;
        RECT 1049.910 2.390 1051.370 4.280 ;
        RECT 1052.210 2.390 1053.670 4.280 ;
        RECT 1054.510 2.390 1055.970 4.280 ;
        RECT 1056.810 2.390 1058.270 4.280 ;
        RECT 1059.110 2.390 1060.570 4.280 ;
        RECT 1061.410 2.390 1062.870 4.280 ;
        RECT 1063.710 2.390 1065.170 4.280 ;
        RECT 1066.010 2.390 1067.470 4.280 ;
        RECT 1068.310 2.390 1069.770 4.280 ;
        RECT 1070.610 2.390 1072.070 4.280 ;
        RECT 1072.910 2.390 1074.370 4.280 ;
        RECT 1075.210 2.390 1076.670 4.280 ;
        RECT 1077.510 2.390 1078.970 4.280 ;
        RECT 1079.810 2.390 1081.270 4.280 ;
        RECT 1082.110 2.390 1083.570 4.280 ;
        RECT 1084.410 2.390 1085.870 4.280 ;
        RECT 1086.710 2.390 1088.170 4.280 ;
        RECT 1089.010 2.390 1090.470 4.280 ;
        RECT 1091.310 2.390 1092.770 4.280 ;
        RECT 1093.610 2.390 1095.070 4.280 ;
        RECT 1095.910 2.390 1097.370 4.280 ;
        RECT 1098.210 2.390 1099.670 4.280 ;
        RECT 1100.510 2.390 1101.970 4.280 ;
        RECT 1102.810 2.390 1104.270 4.280 ;
        RECT 1105.110 2.390 1106.570 4.280 ;
        RECT 1107.410 2.390 1108.870 4.280 ;
        RECT 1109.710 2.390 1111.170 4.280 ;
        RECT 1112.010 2.390 1113.470 4.280 ;
        RECT 1114.310 2.390 1115.770 4.280 ;
        RECT 1116.610 2.390 1118.070 4.280 ;
        RECT 1118.910 2.390 1120.370 4.280 ;
        RECT 1121.210 2.390 1122.670 4.280 ;
        RECT 1123.510 2.390 1124.970 4.280 ;
        RECT 1125.810 2.390 1127.270 4.280 ;
        RECT 1128.110 2.390 1129.570 4.280 ;
        RECT 1130.410 2.390 1131.870 4.280 ;
        RECT 1132.710 2.390 1134.170 4.280 ;
        RECT 1135.010 2.390 1136.470 4.280 ;
        RECT 1137.310 2.390 1138.770 4.280 ;
        RECT 1139.610 2.390 1141.070 4.280 ;
        RECT 1141.910 2.390 1143.370 4.280 ;
        RECT 1144.210 2.390 1145.670 4.280 ;
        RECT 1146.510 2.390 1147.970 4.280 ;
        RECT 1148.810 2.390 1150.270 4.280 ;
        RECT 1151.110 2.390 1152.570 4.280 ;
        RECT 1153.410 2.390 1154.870 4.280 ;
        RECT 1155.710 2.390 1157.170 4.280 ;
        RECT 1158.010 2.390 1159.470 4.280 ;
        RECT 1160.310 2.390 1161.770 4.280 ;
        RECT 1162.610 2.390 1164.070 4.280 ;
        RECT 1164.910 2.390 1166.370 4.280 ;
        RECT 1167.210 2.390 1192.220 4.280 ;
      LAYER met3 ;
        RECT 21.050 4.935 1183.055 1194.585 ;
      LAYER met4 ;
        RECT 80.335 1189.280 1144.185 1194.585 ;
        RECT 80.335 10.240 97.440 1189.280 ;
        RECT 99.840 10.240 174.240 1189.280 ;
        RECT 176.640 10.240 251.040 1189.280 ;
        RECT 253.440 10.240 327.840 1189.280 ;
        RECT 330.240 10.240 404.640 1189.280 ;
        RECT 407.040 10.240 481.440 1189.280 ;
        RECT 483.840 10.240 558.240 1189.280 ;
        RECT 560.640 10.240 635.040 1189.280 ;
        RECT 637.440 10.240 711.840 1189.280 ;
        RECT 714.240 10.240 788.640 1189.280 ;
        RECT 791.040 10.240 865.440 1189.280 ;
        RECT 867.840 10.240 942.240 1189.280 ;
        RECT 944.640 10.240 1019.040 1189.280 ;
        RECT 1021.440 10.240 1095.840 1189.280 ;
        RECT 1098.240 10.240 1144.185 1189.280 ;
        RECT 80.335 4.935 1144.185 10.240 ;
  END
END s3ga_proj
END LIBRARY

