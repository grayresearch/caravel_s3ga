// This is the unpowered netlist.
module x64 (cfg,
    cfgd,
    clk,
    grst,
    io_i,
    io_o,
    rst,
    cfg_i,
    m,
    up_i,
    up_o);
 input cfg;
 output cfgd;
 input clk;
 input grst;
 input io_i;
 output io_o;
 input rst;
 input [4:0] cfg_i;
 input [1:0] m;
 input [15:0] up_i;
 output [7:0] up_o;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire \c.cfg_i_q[0] ;
 wire \c.cfg_i_q[1] ;
 wire \c.cfg_i_q[2] ;
 wire \c.cfg_i_q[3] ;
 wire \c.cfg_i_q[4] ;
 wire \c.genblk1.genblk1.subs.c0.cfg_i_q[0] ;
 wire \c.genblk1.genblk1.subs.c0.cfg_i_q[1] ;
 wire \c.genblk1.genblk1.subs.c0.cfg_i_q[2] ;
 wire \c.genblk1.genblk1.subs.c0.cfg_i_q[3] ;
 wire \c.genblk1.genblk1.subs.c0.cfg_i_q[4] ;
 wire \c.genblk1.genblk1.subs.c0.cfgd ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fd ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fde ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fds ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.m[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.m[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.rst ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fd ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fde ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fds ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fd ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fde ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fds ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fd ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fde ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fds ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.c0.grst ;
 wire \c.genblk1.genblk1.subs.c0.m[0] ;
 wire \c.genblk1.genblk1.subs.c0.m[1] ;
 wire \c.genblk1.genblk1.subs.c0.rst ;
 wire \c.genblk1.genblk1.subs.cs[1].c.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.half_q ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ;
 wire \c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.cfgd ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.o_[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.o_[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.o_[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.o_[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.o_[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.o_[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.o_[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.o_[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.cfgd ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.o_[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.o_[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.o_[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.o_[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.o_[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.o_[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.o_[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.o_[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.cfgd ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.o_[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.o_[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.o_[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.o_[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.o_[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.o_[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.o_[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.o_[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.cfgd ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.o_[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.o_[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.o_[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.o_[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.o_[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.o_[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.o_[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.o_[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[32] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[33] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[34] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[35] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[36] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[37] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[38] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[39] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[9] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o[0] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o[1] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o[2] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o[3] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o[4] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o[5] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o[6] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o[7] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o_[0] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o_[1] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o_[2] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o_[3] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o_[4] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o_[5] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o_[6] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.o_[7] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[0] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[10] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[11] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[14] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[15] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[16] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[17] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[18] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[19] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[1] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[20] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[21] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[22] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[23] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[26] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[27] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[28] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[29] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[2] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[30] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[31] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[3] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[6] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[7] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.o[9] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][0] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][10] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][11] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][12] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][13] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][14] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][15] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][16] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][17] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][18] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][19] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][1] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][20] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][21] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][22] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][23] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][24] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][25] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][26] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][27] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][28] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][29] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][2] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][30] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][31] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][3] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][4] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][5] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][6] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][7] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][8] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][9] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][0] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][10] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][11] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][12] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][13] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][14] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][15] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][16] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][17] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][18] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][19] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][1] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][20] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][21] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][22] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][23] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][24] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][25] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][26] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][27] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][28] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][29] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][2] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][30] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][31] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][3] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][4] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][5] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][6] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][7] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][8] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][9] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][0] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][10] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][11] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][12] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][13] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][14] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][15] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][16] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][17] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][18] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][19] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][1] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][20] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][21] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][22] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][23] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][24] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][25] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][26] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][27] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][28] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][29] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][2] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][30] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][31] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][3] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][4] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][5] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][6] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][7] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][8] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][9] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.seg[0] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.seg[1] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.seg[2] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.seg[4] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[0] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[10] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[11] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[12] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[13] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[14] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[15] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[16] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[17] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[18] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[19] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[1] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[20] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[21] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[22] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[23] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[24] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[25] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[26] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[27] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[28] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[29] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[2] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[30] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[31] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[3] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[4] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[5] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[6] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[7] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[8] ;
 wire \c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[9] ;
 wire clknet_leaf_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_0_1_clk;
 wire clknet_1_1_0_clk;
 wire clknet_1_1_1_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_opt_1_0_clk;
 wire clknet_opt_2_0_clk;
 wire clknet_opt_3_0_clk;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;

 sky130_fd_sc_hd__buf_12 _04814_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[0] ),
    .X(_00170_));
 sky130_fd_sc_hd__buf_8 _04815_ (.A(_00170_),
    .X(_00171_));
 sky130_fd_sc_hd__buf_4 _04816_ (.A(_00171_),
    .X(_00172_));
 sky130_fd_sc_hd__and3b_1 _04817_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[0].x.cfgd ),
    .B(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ),
    .C(\c.genblk1.genblk1.subs.cs[3].c.cfgd ),
    .X(_00173_));
 sky130_fd_sc_hd__clkbuf_2 _04818_ (.A(_00173_),
    .X(_00174_));
 sky130_fd_sc_hd__or2_1 _04819_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[3] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ),
    .X(_00175_));
 sky130_fd_sc_hd__or2_1 _04820_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ),
    .B(_00175_),
    .X(_00176_));
 sky130_fd_sc_hd__or2_1 _04821_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[5] ),
    .B(_00176_),
    .X(_00177_));
 sky130_fd_sc_hd__buf_2 _04822_ (.A(_00177_),
    .X(_00178_));
 sky130_fd_sc_hd__inv_2 _04823_ (.A(_00178_),
    .Y(_00179_));
 sky130_fd_sc_hd__buf_8 _04824_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.rst ),
    .X(_00180_));
 sky130_fd_sc_hd__buf_8 _04825_ (.A(_00180_),
    .X(_00181_));
 sky130_fd_sc_hd__a21o_1 _04826_ (.A1(_00174_),
    .A2(_00179_),
    .B1(_00181_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _04827_ (.A0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[0] ),
    .A1(_00172_),
    .S(_00182_),
    .X(_00183_));
 sky130_fd_sc_hd__clkbuf_1 _04828_ (.A(_00183_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[0] ));
 sky130_fd_sc_hd__buf_6 _04829_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ),
    .X(_00184_));
 sky130_fd_sc_hd__buf_4 _04830_ (.A(_00184_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _04831_ (.A0(net4017),
    .A1(_00185_),
    .S(_00182_),
    .X(_00186_));
 sky130_fd_sc_hd__clkbuf_1 _04832_ (.A(_00186_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[1] ));
 sky130_fd_sc_hd__buf_12 _04833_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[2] ),
    .X(_00187_));
 sky130_fd_sc_hd__buf_6 _04834_ (.A(_00187_),
    .X(_00188_));
 sky130_fd_sc_hd__buf_4 _04835_ (.A(_00188_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _04836_ (.A0(net3672),
    .A1(_00189_),
    .S(_00182_),
    .X(_00190_));
 sky130_fd_sc_hd__clkbuf_1 _04837_ (.A(_00190_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[2] ));
 sky130_fd_sc_hd__buf_6 _04838_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ),
    .X(_00191_));
 sky130_fd_sc_hd__clkbuf_4 _04839_ (.A(_00191_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _04840_ (.A0(net4021),
    .A1(_00192_),
    .S(_00182_),
    .X(_00193_));
 sky130_fd_sc_hd__clkbuf_1 _04841_ (.A(_00193_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[3] ));
 sky130_fd_sc_hd__inv_2 _04842_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.rst ),
    .Y(_00194_));
 sky130_fd_sc_hd__buf_4 _04843_ (.A(_00194_),
    .X(_00195_));
 sky130_fd_sc_hd__buf_6 _04844_ (.A(_00195_),
    .X(_00196_));
 sky130_fd_sc_hd__buf_2 _04845_ (.A(_00196_),
    .X(_00197_));
 sky130_fd_sc_hd__clkbuf_2 _04846_ (.A(net3786),
    .X(_00198_));
 sky130_fd_sc_hd__nor3b_2 _04847_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ),
    .B(_00198_),
    .C_N(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ),
    .Y(_00199_));
 sky130_fd_sc_hd__nand2_1 _04848_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[5] ),
    .B(_00176_),
    .Y(_00200_));
 sky130_fd_sc_hd__and3_2 _04849_ (.A(_00174_),
    .B(_00178_),
    .C(_00200_),
    .X(_00201_));
 sky130_fd_sc_hd__nand2_2 _04850_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[0] ),
    .B(_00178_),
    .Y(_00202_));
 sky130_fd_sc_hd__inv_2 _04851_ (.A(_00202_),
    .Y(_00203_));
 sky130_fd_sc_hd__or3b_2 _04852_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ),
    .B(_00198_),
    .C_N(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ),
    .X(_00204_));
 sky130_fd_sc_hd__or3b_2 _04853_ (.A(_00204_),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[5] ),
    .C_N(_00174_),
    .X(_00205_));
 sky130_fd_sc_hd__a32o_1 _04854_ (.A1(_00199_),
    .A2(_00201_),
    .A3(_00203_),
    .B1(_00205_),
    .B2(net3415),
    .X(_00206_));
 sky130_fd_sc_hd__and2_1 _04855_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[0] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.rst ),
    .X(_00207_));
 sky130_fd_sc_hd__clkbuf_2 _04856_ (.A(_00207_),
    .X(_00208_));
 sky130_fd_sc_hd__buf_4 _04857_ (.A(_00208_),
    .X(_00209_));
 sky130_fd_sc_hd__buf_8 _04858_ (.A(_00209_),
    .X(_00210_));
 sky130_fd_sc_hd__a21o_1 _04859_ (.A1(_00197_),
    .A2(_00206_),
    .B1(_00210_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[4] ));
 sky130_fd_sc_hd__buf_12 _04860_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ),
    .X(_00211_));
 sky130_fd_sc_hd__and2_1 _04861_ (.A(_00211_),
    .B(_00178_),
    .X(_00212_));
 sky130_fd_sc_hd__a32o_1 _04862_ (.A1(_00199_),
    .A2(_00201_),
    .A3(_00212_),
    .B1(_00205_),
    .B2(net4174),
    .X(_00213_));
 sky130_fd_sc_hd__and2_1 _04863_ (.A(_00180_),
    .B(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ),
    .X(_00214_));
 sky130_fd_sc_hd__clkbuf_4 _04864_ (.A(_00214_),
    .X(_00215_));
 sky130_fd_sc_hd__clkbuf_8 _04865_ (.A(_00215_),
    .X(_00216_));
 sky130_fd_sc_hd__a21o_1 _04866_ (.A1(_00197_),
    .A2(_00213_),
    .B1(_00216_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[5] ));
 sky130_fd_sc_hd__nand2_2 _04867_ (.A(net3667),
    .B(_00178_),
    .Y(_00217_));
 sky130_fd_sc_hd__inv_2 _04868_ (.A(_00217_),
    .Y(_00218_));
 sky130_fd_sc_hd__a32o_1 _04869_ (.A1(_00199_),
    .A2(_00201_),
    .A3(_00218_),
    .B1(_00205_),
    .B2(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ),
    .X(_00219_));
 sky130_fd_sc_hd__and2_1 _04870_ (.A(_00180_),
    .B(\c.genblk1.genblk1.subs.c0.cfg_i_q[2] ),
    .X(_00220_));
 sky130_fd_sc_hd__buf_4 _04871_ (.A(_00220_),
    .X(_00221_));
 sky130_fd_sc_hd__buf_4 _04872_ (.A(_00221_),
    .X(_00222_));
 sky130_fd_sc_hd__a21o_1 _04873_ (.A1(_00197_),
    .A2(_00219_),
    .B1(_00222_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[6] ));
 sky130_fd_sc_hd__clkbuf_4 _04874_ (.A(_00195_),
    .X(_00223_));
 sky130_fd_sc_hd__and2_1 _04875_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ),
    .B(_00178_),
    .X(_00224_));
 sky130_fd_sc_hd__a32o_1 _04876_ (.A1(_00199_),
    .A2(_00201_),
    .A3(_00224_),
    .B1(_00205_),
    .B2(net4157),
    .X(_00225_));
 sky130_fd_sc_hd__nand2_4 _04877_ (.A(_00180_),
    .B(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ),
    .Y(_00226_));
 sky130_fd_sc_hd__buf_4 _04878_ (.A(_00226_),
    .X(_00227_));
 sky130_fd_sc_hd__a21bo_1 _04879_ (.A1(_00223_),
    .A2(_00225_),
    .B1_N(_00227_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[7] ));
 sky130_fd_sc_hd__buf_6 _04880_ (.A(_00181_),
    .X(_00228_));
 sky130_fd_sc_hd__buf_4 _04881_ (.A(_00228_),
    .X(_00229_));
 sky130_fd_sc_hd__inv_2 _04882_ (.A(net3998),
    .Y(_00230_));
 sky130_fd_sc_hd__and2_1 _04883_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ),
    .B(_00175_),
    .X(_00231_));
 sky130_fd_sc_hd__or4bb_2 _04884_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[5] ),
    .B(_00231_),
    .C_N(_00174_),
    .D_N(_00176_),
    .X(_00232_));
 sky130_fd_sc_hd__or3b_4 _04885_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ),
    .B(_00232_),
    .C_N(_00198_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _04886_ (.A0(_00202_),
    .A1(_00230_),
    .S(_00233_),
    .X(_00234_));
 sky130_fd_sc_hd__buf_8 _04887_ (.A(_00170_),
    .X(_00235_));
 sky130_fd_sc_hd__buf_12 _04888_ (.A(_00180_),
    .X(_00236_));
 sky130_fd_sc_hd__nand2_8 _04889_ (.A(_00235_),
    .B(_00236_),
    .Y(_00237_));
 sky130_fd_sc_hd__clkbuf_4 _04890_ (.A(_00237_),
    .X(_00238_));
 sky130_fd_sc_hd__o21ai_1 _04891_ (.A1(_00229_),
    .A2(_00234_),
    .B1(_00238_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[8] ));
 sky130_fd_sc_hd__mux2_1 _04892_ (.A0(_00212_),
    .A1(net4213),
    .S(_00233_),
    .X(_00239_));
 sky130_fd_sc_hd__a21o_1 _04893_ (.A1(_00197_),
    .A2(_00239_),
    .B1(_00216_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[9] ));
 sky130_fd_sc_hd__mux2_1 _04894_ (.A0(_00218_),
    .A1(net4178),
    .S(_00233_),
    .X(_00240_));
 sky130_fd_sc_hd__a21o_1 _04895_ (.A1(_00197_),
    .A2(_00240_),
    .B1(_00222_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[10] ));
 sky130_fd_sc_hd__mux2_1 _04896_ (.A0(_00224_),
    .A1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ),
    .S(_00233_),
    .X(_00241_));
 sky130_fd_sc_hd__a21bo_1 _04897_ (.A1(_00223_),
    .A2(_00241_),
    .B1_N(_00227_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[11] ));
 sky130_fd_sc_hd__inv_2 _04898_ (.A(net3896),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _04899_ (.A(_00198_),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ),
    .Y(_00243_));
 sky130_fd_sc_hd__nor2_2 _04900_ (.A(_00232_),
    .B(_00243_),
    .Y(_00244_));
 sky130_fd_sc_hd__mux2_1 _04901_ (.A0(_00242_),
    .A1(_00202_),
    .S(_00244_),
    .X(_00245_));
 sky130_fd_sc_hd__o21ai_1 _04902_ (.A1(_00229_),
    .A2(_00245_),
    .B1(_00238_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _04903_ (.A0(net4197),
    .A1(_00212_),
    .S(_00244_),
    .X(_00246_));
 sky130_fd_sc_hd__a21o_1 _04904_ (.A1(_00197_),
    .A2(_00246_),
    .B1(_00216_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[13] ));
 sky130_fd_sc_hd__inv_2 _04905_ (.A(net3663),
    .Y(_00247_));
 sky130_fd_sc_hd__mux2_1 _04906_ (.A0(_00247_),
    .A1(_00217_),
    .S(_00244_),
    .X(_00248_));
 sky130_fd_sc_hd__buf_4 _04907_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.rst ),
    .X(_00249_));
 sky130_fd_sc_hd__nand2_1 _04908_ (.A(_00249_),
    .B(_00187_),
    .Y(_00250_));
 sky130_fd_sc_hd__buf_6 _04909_ (.A(_00250_),
    .X(_00251_));
 sky130_fd_sc_hd__buf_4 _04910_ (.A(_00251_),
    .X(_00252_));
 sky130_fd_sc_hd__o21ai_1 _04911_ (.A1(_00229_),
    .A2(_00248_),
    .B1(_00252_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _04912_ (.A0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ),
    .A1(_00224_),
    .S(_00244_),
    .X(_00253_));
 sky130_fd_sc_hd__a21bo_1 _04913_ (.A1(_00223_),
    .A2(_00253_),
    .B1_N(_00227_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[15] ));
 sky130_fd_sc_hd__nor2_2 _04914_ (.A(_00175_),
    .B(_00232_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _04915_ (.A(_00202_),
    .B(_00254_),
    .Y(_00255_));
 sky130_fd_sc_hd__or2_1 _04916_ (.A(net4072),
    .B(_00254_),
    .X(_00256_));
 sky130_fd_sc_hd__a31o_1 _04917_ (.A1(_00223_),
    .A2(_00255_),
    .A3(_00256_),
    .B1(_00210_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _04918_ (.A(_00184_),
    .B(_00178_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand2_1 _04919_ (.A(_00257_),
    .B(_00254_),
    .Y(_00258_));
 sky130_fd_sc_hd__or2_1 _04920_ (.A(net4063),
    .B(_00254_),
    .X(_00259_));
 sky130_fd_sc_hd__a31o_1 _04921_ (.A1(_00223_),
    .A2(_00258_),
    .A3(_00259_),
    .B1(_00216_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _04922_ (.A(_00217_),
    .B(_00254_),
    .Y(_00260_));
 sky130_fd_sc_hd__or2_1 _04923_ (.A(net4176),
    .B(_00254_),
    .X(_00261_));
 sky130_fd_sc_hd__buf_6 _04924_ (.A(_00221_),
    .X(_00262_));
 sky130_fd_sc_hd__a31o_1 _04925_ (.A1(_00223_),
    .A2(_00260_),
    .A3(_00261_),
    .B1(_00262_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[18] ));
 sky130_fd_sc_hd__buf_6 _04926_ (.A(_00227_),
    .X(_00263_));
 sky130_fd_sc_hd__buf_12 _04927_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ),
    .X(_00264_));
 sky130_fd_sc_hd__nand2_1 _04928_ (.A(_00264_),
    .B(_00178_),
    .Y(_00265_));
 sky130_fd_sc_hd__nor2_1 _04929_ (.A(net3725),
    .B(_00254_),
    .Y(_00266_));
 sky130_fd_sc_hd__buf_12 _04930_ (.A(_00180_),
    .X(_00267_));
 sky130_fd_sc_hd__buf_6 _04931_ (.A(_00267_),
    .X(_00268_));
 sky130_fd_sc_hd__a211o_1 _04932_ (.A1(_00265_),
    .A2(_00254_),
    .B1(_00266_),
    .C1(_00268_),
    .X(_00269_));
 sky130_fd_sc_hd__nand2_1 _04933_ (.A(_00263_),
    .B(_00269_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[19] ));
 sky130_fd_sc_hd__and4b_2 _04934_ (.A_N(_00198_),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ),
    .C(_00201_),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _04935_ (.A0(net4148),
    .A1(_00203_),
    .S(_00270_),
    .X(_00271_));
 sky130_fd_sc_hd__a21o_1 _04936_ (.A1(_00197_),
    .A2(_00271_),
    .B1(_00210_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _04937_ (.A0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ),
    .A1(_00212_),
    .S(_00270_),
    .X(_00272_));
 sky130_fd_sc_hd__a21o_1 _04938_ (.A1(_00197_),
    .A2(_00272_),
    .B1(_00216_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _04939_ (.A0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ),
    .A1(_00218_),
    .S(_00270_),
    .X(_00273_));
 sky130_fd_sc_hd__a21o_1 _04940_ (.A1(_00197_),
    .A2(_00273_),
    .B1(_00222_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[22] ));
 sky130_fd_sc_hd__inv_2 _04941_ (.A(net3787),
    .Y(_00274_));
 sky130_fd_sc_hd__mux2_1 _04942_ (.A0(_00274_),
    .A1(_00265_),
    .S(_00270_),
    .X(_00275_));
 sky130_fd_sc_hd__buf_4 _04943_ (.A(_00226_),
    .X(_00276_));
 sky130_fd_sc_hd__o21ai_1 _04944_ (.A1(_00229_),
    .A2(_00275_),
    .B1(_00276_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4b_2 _04945_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ),
    .B(_00201_),
    .C(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ),
    .D(_00198_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _04946_ (.A0(net3390),
    .A1(_00203_),
    .S(_00277_),
    .X(_00278_));
 sky130_fd_sc_hd__a21o_1 _04947_ (.A1(_00197_),
    .A2(_00278_),
    .B1(_00210_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[24] ));
 sky130_fd_sc_hd__buf_4 _04948_ (.A(_00196_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _04949_ (.A0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ),
    .A1(_00212_),
    .S(_00277_),
    .X(_00280_));
 sky130_fd_sc_hd__a21o_1 _04950_ (.A1(_00279_),
    .A2(_00280_),
    .B1(_00216_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _04951_ (.A0(net4200),
    .A1(_00218_),
    .S(_00277_),
    .X(_00281_));
 sky130_fd_sc_hd__a21o_1 _04952_ (.A1(_00279_),
    .A2(_00281_),
    .B1(_00222_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _04953_ (.A0(net4038),
    .A1(_00224_),
    .S(_00277_),
    .X(_00282_));
 sky130_fd_sc_hd__a21bo_1 _04954_ (.A1(_00223_),
    .A2(_00282_),
    .B1_N(_00227_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[27] ));
 sky130_fd_sc_hd__and4_2 _04955_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ),
    .B(_00198_),
    .C(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ),
    .D(_00201_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _04956_ (.A0(net4139),
    .A1(_00203_),
    .S(_00283_),
    .X(_00284_));
 sky130_fd_sc_hd__a21o_1 _04957_ (.A1(_00279_),
    .A2(_00284_),
    .B1(_00210_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _04958_ (.A0(net3494),
    .A1(_00212_),
    .S(_00283_),
    .X(_00285_));
 sky130_fd_sc_hd__a21o_1 _04959_ (.A1(_00279_),
    .A2(_00285_),
    .B1(_00216_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _04960_ (.A0(net4122),
    .A1(_00218_),
    .S(_00283_),
    .X(_00286_));
 sky130_fd_sc_hd__a21o_1 _04961_ (.A1(_00279_),
    .A2(_00286_),
    .B1(_00222_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _04962_ (.A0(net4094),
    .A1(_00224_),
    .S(_00283_),
    .X(_00287_));
 sky130_fd_sc_hd__a21bo_1 _04963_ (.A1(_00223_),
    .A2(_00287_),
    .B1_N(_00227_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[31] ));
 sky130_fd_sc_hd__buf_4 _04964_ (.A(_00235_),
    .X(_00288_));
 sky130_fd_sc_hd__nand2_1 _04965_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[5] ),
    .B(_00174_),
    .Y(_00289_));
 sky130_fd_sc_hd__o21a_2 _04966_ (.A1(_00176_),
    .A2(_00289_),
    .B1(_00195_),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _04967_ (.A0(_00288_),
    .A1(net3788),
    .S(_00290_),
    .X(_00291_));
 sky130_fd_sc_hd__clkbuf_1 _04968_ (.A(_00291_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[32] ));
 sky130_fd_sc_hd__buf_8 _04969_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ),
    .X(_00292_));
 sky130_fd_sc_hd__buf_4 _04970_ (.A(_00292_),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _04971_ (.A0(_00293_),
    .A1(net4051),
    .S(_00290_),
    .X(_00294_));
 sky130_fd_sc_hd__clkbuf_1 _04972_ (.A(_00294_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[33] ));
 sky130_fd_sc_hd__buf_4 _04973_ (.A(_00188_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _04974_ (.A0(_00295_),
    .A1(net3764),
    .S(_00290_),
    .X(_00296_));
 sky130_fd_sc_hd__clkbuf_1 _04975_ (.A(_00296_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[34] ));
 sky130_fd_sc_hd__buf_6 _04976_ (.A(_00191_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _04977_ (.A0(_00297_),
    .A1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[35] ),
    .S(_00290_),
    .X(_00298_));
 sky130_fd_sc_hd__clkbuf_1 _04978_ (.A(_00298_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[35] ));
 sky130_fd_sc_hd__a21bo_1 _04979_ (.A1(_00178_),
    .A2(_00200_),
    .B1_N(_00174_),
    .X(_00299_));
 sky130_fd_sc_hd__nor2_1 _04980_ (.A(_00204_),
    .B(_00289_),
    .Y(_00300_));
 sky130_fd_sc_hd__inv_2 _04981_ (.A(net3977),
    .Y(_00301_));
 sky130_fd_sc_hd__o32a_1 _04982_ (.A1(_00204_),
    .A2(_00202_),
    .A3(_00299_),
    .B1(_00300_),
    .B2(_00301_),
    .X(_00302_));
 sky130_fd_sc_hd__o21ai_1 _04983_ (.A1(_00229_),
    .A2(_00302_),
    .B1(_00238_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[36] ));
 sky130_fd_sc_hd__inv_2 _04984_ (.A(net3818),
    .Y(_00303_));
 sky130_fd_sc_hd__o32a_1 _04985_ (.A1(_00204_),
    .A2(_00257_),
    .A3(_00299_),
    .B1(_00300_),
    .B2(_00303_),
    .X(_00304_));
 sky130_fd_sc_hd__nand2_8 _04986_ (.A(_00236_),
    .B(_00292_),
    .Y(_00305_));
 sky130_fd_sc_hd__clkbuf_4 _04987_ (.A(_00305_),
    .X(_00306_));
 sky130_fd_sc_hd__o21ai_1 _04988_ (.A1(_00229_),
    .A2(_00304_),
    .B1(_00306_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[37] ));
 sky130_fd_sc_hd__inv_2 _04989_ (.A(net4012),
    .Y(_00307_));
 sky130_fd_sc_hd__o32a_1 _04990_ (.A1(_00204_),
    .A2(_00217_),
    .A3(_00299_),
    .B1(_00300_),
    .B2(_00307_),
    .X(_00308_));
 sky130_fd_sc_hd__o21ai_1 _04991_ (.A1(_00229_),
    .A2(_00308_),
    .B1(_00252_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[38] ));
 sky130_fd_sc_hd__inv_2 _04992_ (.A(net3631),
    .Y(_00309_));
 sky130_fd_sc_hd__o32a_1 _04993_ (.A1(_00204_),
    .A2(_00265_),
    .A3(_00299_),
    .B1(_00300_),
    .B2(_00309_),
    .X(_00310_));
 sky130_fd_sc_hd__o21ai_1 _04994_ (.A1(_00229_),
    .A2(_00310_),
    .B1(_00276_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[39] ));
 sky130_fd_sc_hd__clkbuf_16 _04995_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ),
    .X(_00311_));
 sky130_fd_sc_hd__and3b_1 _04996_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[1].x.cfgd ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.cfgd ),
    .C(_00311_),
    .X(_00312_));
 sky130_fd_sc_hd__buf_2 _04997_ (.A(_00312_),
    .X(_00313_));
 sky130_fd_sc_hd__or2_1 _04998_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ),
    .X(_00314_));
 sky130_fd_sc_hd__or2_1 _04999_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[4] ),
    .B(_00314_),
    .X(_00315_));
 sky130_fd_sc_hd__or2_1 _05000_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[5] ),
    .B(_00315_),
    .X(_00316_));
 sky130_fd_sc_hd__clkbuf_4 _05001_ (.A(_00316_),
    .X(_00317_));
 sky130_fd_sc_hd__inv_2 _05002_ (.A(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__a21oi_4 _05003_ (.A1(_00313_),
    .A2(_00318_),
    .B1(_00267_),
    .Y(_00319_));
 sky130_fd_sc_hd__mux2_1 _05004_ (.A0(_00288_),
    .A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[0] ),
    .S(_00319_),
    .X(_00320_));
 sky130_fd_sc_hd__clkbuf_1 _05005_ (.A(_00320_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _05006_ (.A0(_00293_),
    .A1(net4018),
    .S(_00319_),
    .X(_00321_));
 sky130_fd_sc_hd__clkbuf_1 _05007_ (.A(_00321_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _05008_ (.A0(_00295_),
    .A1(net3964),
    .S(_00319_),
    .X(_00322_));
 sky130_fd_sc_hd__clkbuf_1 _05009_ (.A(_00322_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _05010_ (.A0(_00297_),
    .A1(net4124),
    .S(_00319_),
    .X(_00323_));
 sky130_fd_sc_hd__clkbuf_1 _05011_ (.A(_00323_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[3] ));
 sky130_fd_sc_hd__or3b_1 _05012_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[4] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ),
    .C_N(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ),
    .X(_00324_));
 sky130_fd_sc_hd__buf_2 _05013_ (.A(_00324_),
    .X(_00325_));
 sky130_fd_sc_hd__nand2_1 _05014_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[5] ),
    .B(_00315_),
    .Y(_00326_));
 sky130_fd_sc_hd__and2_1 _05015_ (.A(_00317_),
    .B(_00326_),
    .X(_00327_));
 sky130_fd_sc_hd__nand2_1 _05016_ (.A(_00313_),
    .B(_00327_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_2 _05017_ (.A(_00170_),
    .B(_00317_),
    .Y(_00329_));
 sky130_fd_sc_hd__inv_2 _05018_ (.A(_00325_),
    .Y(_00330_));
 sky130_fd_sc_hd__and3b_1 _05019_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[5] ),
    .B(_00313_),
    .C(_00330_),
    .X(_00331_));
 sky130_fd_sc_hd__inv_2 _05020_ (.A(net3554),
    .Y(_00332_));
 sky130_fd_sc_hd__o32a_1 _05021_ (.A1(_00325_),
    .A2(_00328_),
    .A3(_00329_),
    .B1(_00331_),
    .B2(_00332_),
    .X(_00333_));
 sky130_fd_sc_hd__o21ai_1 _05022_ (.A1(_00229_),
    .A2(_00333_),
    .B1(_00238_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[4] ));
 sky130_fd_sc_hd__buf_2 _05023_ (.A(_00228_),
    .X(_00334_));
 sky130_fd_sc_hd__nand2_4 _05024_ (.A(_00211_),
    .B(_00317_),
    .Y(_00335_));
 sky130_fd_sc_hd__inv_2 _05025_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ),
    .Y(_00336_));
 sky130_fd_sc_hd__o32a_1 _05026_ (.A1(_00325_),
    .A2(_00328_),
    .A3(_00335_),
    .B1(_00331_),
    .B2(_00336_),
    .X(_00337_));
 sky130_fd_sc_hd__o21ai_1 _05027_ (.A1(_00334_),
    .A2(_00337_),
    .B1(_00306_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[5] ));
 sky130_fd_sc_hd__nand2_2 _05028_ (.A(_00187_),
    .B(_00317_),
    .Y(_00338_));
 sky130_fd_sc_hd__inv_2 _05029_ (.A(net4131),
    .Y(_00339_));
 sky130_fd_sc_hd__o32a_1 _05030_ (.A1(_00325_),
    .A2(_00328_),
    .A3(_00338_),
    .B1(_00331_),
    .B2(_00339_),
    .X(_00340_));
 sky130_fd_sc_hd__o21ai_1 _05031_ (.A1(_00334_),
    .A2(_00340_),
    .B1(_00252_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[6] ));
 sky130_fd_sc_hd__nand2_2 _05032_ (.A(_00264_),
    .B(_00317_),
    .Y(_00341_));
 sky130_fd_sc_hd__inv_2 _05033_ (.A(net4136),
    .Y(_00342_));
 sky130_fd_sc_hd__o32a_1 _05034_ (.A1(_00325_),
    .A2(_00328_),
    .A3(_00341_),
    .B1(_00331_),
    .B2(_00342_),
    .X(_00343_));
 sky130_fd_sc_hd__o21ai_1 _05035_ (.A1(_00334_),
    .A2(_00343_),
    .B1(_00276_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _05036_ (.A(net3945),
    .Y(_00344_));
 sky130_fd_sc_hd__and2_1 _05037_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[4] ),
    .B(_00314_),
    .X(_00345_));
 sky130_fd_sc_hd__or4bb_2 _05038_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[5] ),
    .B(_00345_),
    .C_N(_00312_),
    .D_N(_00315_),
    .X(_00346_));
 sky130_fd_sc_hd__or3b_2 _05039_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ),
    .B(_00346_),
    .C_N(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _05040_ (.A0(_00329_),
    .A1(_00344_),
    .S(_00347_),
    .X(_00348_));
 sky130_fd_sc_hd__o21ai_1 _05041_ (.A1(_00334_),
    .A2(_00348_),
    .B1(_00238_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[8] ));
 sky130_fd_sc_hd__inv_2 _05042_ (.A(net3618),
    .Y(_00349_));
 sky130_fd_sc_hd__mux2_1 _05043_ (.A0(_00335_),
    .A1(_00349_),
    .S(_00347_),
    .X(_00350_));
 sky130_fd_sc_hd__o21ai_1 _05044_ (.A1(_00334_),
    .A2(_00350_),
    .B1(_00306_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[9] ));
 sky130_fd_sc_hd__inv_2 _05045_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ),
    .Y(_00351_));
 sky130_fd_sc_hd__mux2_1 _05046_ (.A0(_00338_),
    .A1(_00351_),
    .S(_00347_),
    .X(_00352_));
 sky130_fd_sc_hd__o21ai_1 _05047_ (.A1(_00334_),
    .A2(_00352_),
    .B1(_00252_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[10] ));
 sky130_fd_sc_hd__clkinv_2 _05048_ (.A(net4118),
    .Y(_00353_));
 sky130_fd_sc_hd__mux2_1 _05049_ (.A0(_00341_),
    .A1(_00353_),
    .S(_00347_),
    .X(_00354_));
 sky130_fd_sc_hd__o21ai_1 _05050_ (.A1(_00334_),
    .A2(_00354_),
    .B1(_00276_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[11] ));
 sky130_fd_sc_hd__inv_2 _05051_ (.A(net3245),
    .Y(_00355_));
 sky130_fd_sc_hd__nand2_1 _05052_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ),
    .Y(_00356_));
 sky130_fd_sc_hd__nor2_2 _05053_ (.A(_00346_),
    .B(_00356_),
    .Y(_00357_));
 sky130_fd_sc_hd__mux2_1 _05054_ (.A0(_00355_),
    .A1(_00329_),
    .S(_00357_),
    .X(_00358_));
 sky130_fd_sc_hd__o21ai_1 _05055_ (.A1(_00334_),
    .A2(_00358_),
    .B1(_00238_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[12] ));
 sky130_fd_sc_hd__inv_2 _05056_ (.A(net3341),
    .Y(_00359_));
 sky130_fd_sc_hd__mux2_1 _05057_ (.A0(_00359_),
    .A1(_00335_),
    .S(_00357_),
    .X(_00360_));
 sky130_fd_sc_hd__o21ai_1 _05058_ (.A1(_00334_),
    .A2(_00360_),
    .B1(_00306_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[13] ));
 sky130_fd_sc_hd__inv_2 _05059_ (.A(net3168),
    .Y(_00361_));
 sky130_fd_sc_hd__mux2_1 _05060_ (.A0(_00361_),
    .A1(_00338_),
    .S(_00357_),
    .X(_00362_));
 sky130_fd_sc_hd__o21ai_1 _05061_ (.A1(_00334_),
    .A2(_00362_),
    .B1(_00252_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[14] ));
 sky130_fd_sc_hd__buf_6 _05062_ (.A(_00181_),
    .X(_00363_));
 sky130_fd_sc_hd__buf_2 _05063_ (.A(_00363_),
    .X(_00364_));
 sky130_fd_sc_hd__inv_2 _05064_ (.A(net4185),
    .Y(_00365_));
 sky130_fd_sc_hd__mux2_1 _05065_ (.A0(_00365_),
    .A1(_00341_),
    .S(_00357_),
    .X(_00366_));
 sky130_fd_sc_hd__o21ai_1 _05066_ (.A1(_00364_),
    .A2(_00366_),
    .B1(_00276_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[15] ));
 sky130_fd_sc_hd__buf_4 _05067_ (.A(_00196_),
    .X(_00367_));
 sky130_fd_sc_hd__nor2_2 _05068_ (.A(_00314_),
    .B(_00346_),
    .Y(_00368_));
 sky130_fd_sc_hd__nand2_1 _05069_ (.A(_00329_),
    .B(_00368_),
    .Y(_00369_));
 sky130_fd_sc_hd__or2_1 _05070_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ),
    .B(_00368_),
    .X(_00370_));
 sky130_fd_sc_hd__a31o_1 _05071_ (.A1(_00367_),
    .A2(_00369_),
    .A3(_00370_),
    .B1(_00210_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _05072_ (.A(_00335_),
    .B(_00368_),
    .Y(_00371_));
 sky130_fd_sc_hd__or2_1 _05073_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[17] ),
    .B(_00368_),
    .X(_00372_));
 sky130_fd_sc_hd__a31o_1 _05074_ (.A1(_00367_),
    .A2(_00371_),
    .A3(_00372_),
    .B1(_00216_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _05075_ (.A(_00338_),
    .B(_00368_),
    .Y(_00373_));
 sky130_fd_sc_hd__or2_1 _05076_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[18] ),
    .B(_00368_),
    .X(_00374_));
 sky130_fd_sc_hd__a31o_1 _05077_ (.A1(_00367_),
    .A2(_00373_),
    .A3(_00374_),
    .B1(_00262_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _05078_ (.A(net3677),
    .B(_00368_),
    .Y(_00375_));
 sky130_fd_sc_hd__a211o_1 _05079_ (.A1(_00341_),
    .A2(_00368_),
    .B1(_00375_),
    .C1(_00268_),
    .X(_00376_));
 sky130_fd_sc_hd__nand2_1 _05080_ (.A(_00263_),
    .B(_00376_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[19] ));
 sky130_fd_sc_hd__inv_2 _05081_ (.A(net4079),
    .Y(_00377_));
 sky130_fd_sc_hd__and3_1 _05082_ (.A(_00313_),
    .B(_00317_),
    .C(_00326_),
    .X(_00378_));
 sky130_fd_sc_hd__and4b_1 _05083_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ),
    .C(_00378_),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[4] ),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _05084_ (.A0(_00377_),
    .A1(_00329_),
    .S(_00379_),
    .X(_00380_));
 sky130_fd_sc_hd__o21ai_1 _05085_ (.A1(_00364_),
    .A2(_00380_),
    .B1(_00238_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[20] ));
 sky130_fd_sc_hd__or2_1 _05086_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ),
    .B(_00379_),
    .X(_00381_));
 sky130_fd_sc_hd__nand2_1 _05087_ (.A(_00335_),
    .B(_00379_),
    .Y(_00382_));
 sky130_fd_sc_hd__a31o_1 _05088_ (.A1(_00367_),
    .A2(_00381_),
    .A3(_00382_),
    .B1(_00216_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[21] ));
 sky130_fd_sc_hd__inv_2 _05089_ (.A(net3995),
    .Y(_00383_));
 sky130_fd_sc_hd__mux2_1 _05090_ (.A0(_00383_),
    .A1(_00338_),
    .S(_00379_),
    .X(_00384_));
 sky130_fd_sc_hd__o21ai_1 _05091_ (.A1(_00364_),
    .A2(_00384_),
    .B1(_00252_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[22] ));
 sky130_fd_sc_hd__inv_2 _05092_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[23] ),
    .Y(_00385_));
 sky130_fd_sc_hd__mux2_1 _05093_ (.A0(_00385_),
    .A1(_00341_),
    .S(_00379_),
    .X(_00386_));
 sky130_fd_sc_hd__o21ai_1 _05094_ (.A1(_00364_),
    .A2(_00386_),
    .B1(_00276_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[23] ));
 sky130_fd_sc_hd__inv_2 _05095_ (.A(net3700),
    .Y(_00387_));
 sky130_fd_sc_hd__and4b_2 _05096_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ),
    .B(_00378_),
    .C(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[4] ),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _05097_ (.A0(_00387_),
    .A1(_00329_),
    .S(_00388_),
    .X(_00389_));
 sky130_fd_sc_hd__o21ai_1 _05098_ (.A1(_00364_),
    .A2(_00389_),
    .B1(_00238_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[24] ));
 sky130_fd_sc_hd__inv_2 _05099_ (.A(net4114),
    .Y(_00390_));
 sky130_fd_sc_hd__mux2_1 _05100_ (.A0(_00390_),
    .A1(_00335_),
    .S(_00388_),
    .X(_00391_));
 sky130_fd_sc_hd__o21ai_1 _05101_ (.A1(_00364_),
    .A2(_00391_),
    .B1(_00306_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[25] ));
 sky130_fd_sc_hd__nand2_1 _05102_ (.A(_00338_),
    .B(_00388_),
    .Y(_00392_));
 sky130_fd_sc_hd__or2_1 _05103_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ),
    .B(_00388_),
    .X(_00393_));
 sky130_fd_sc_hd__buf_8 _05104_ (.A(_00221_),
    .X(_00394_));
 sky130_fd_sc_hd__a31o_1 _05105_ (.A1(_00367_),
    .A2(_00392_),
    .A3(_00393_),
    .B1(_00394_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[26] ));
 sky130_fd_sc_hd__inv_2 _05106_ (.A(net4099),
    .Y(_00395_));
 sky130_fd_sc_hd__mux2_1 _05107_ (.A0(_00395_),
    .A1(_00341_),
    .S(_00388_),
    .X(_00396_));
 sky130_fd_sc_hd__o21ai_1 _05108_ (.A1(_00364_),
    .A2(_00396_),
    .B1(_00276_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[27] ));
 sky130_fd_sc_hd__inv_2 _05109_ (.A(net4209),
    .Y(_00397_));
 sky130_fd_sc_hd__and4_2 _05110_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[4] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ),
    .C(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ),
    .D(_00378_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _05111_ (.A0(_00397_),
    .A1(_00329_),
    .S(_00398_),
    .X(_00399_));
 sky130_fd_sc_hd__o21ai_1 _05112_ (.A1(_00364_),
    .A2(_00399_),
    .B1(_00238_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[28] ));
 sky130_fd_sc_hd__inv_2 _05113_ (.A(net3575),
    .Y(_00400_));
 sky130_fd_sc_hd__mux2_1 _05114_ (.A0(_00400_),
    .A1(_00335_),
    .S(_00398_),
    .X(_00401_));
 sky130_fd_sc_hd__o21ai_1 _05115_ (.A1(_00364_),
    .A2(_00401_),
    .B1(_00306_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[29] ));
 sky130_fd_sc_hd__inv_2 _05116_ (.A(net4138),
    .Y(_00402_));
 sky130_fd_sc_hd__mux2_1 _05117_ (.A0(_00402_),
    .A1(_00338_),
    .S(_00398_),
    .X(_00403_));
 sky130_fd_sc_hd__o21ai_1 _05118_ (.A1(_00364_),
    .A2(_00403_),
    .B1(_00252_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[30] ));
 sky130_fd_sc_hd__nor2_1 _05119_ (.A(net4158),
    .B(_00398_),
    .Y(_00404_));
 sky130_fd_sc_hd__a211o_1 _05120_ (.A1(_00341_),
    .A2(_00398_),
    .B1(_00404_),
    .C1(_00268_),
    .X(_00405_));
 sky130_fd_sc_hd__nand2_1 _05121_ (.A(_00263_),
    .B(_00405_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[31] ));
 sky130_fd_sc_hd__nand2_1 _05122_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[5] ),
    .B(_00313_),
    .Y(_00406_));
 sky130_fd_sc_hd__buf_6 _05123_ (.A(_00194_),
    .X(_00407_));
 sky130_fd_sc_hd__buf_6 _05124_ (.A(_00407_),
    .X(_00408_));
 sky130_fd_sc_hd__o21a_2 _05125_ (.A1(_00315_),
    .A2(_00406_),
    .B1(_00408_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _05126_ (.A0(_00288_),
    .A1(net4078),
    .S(_00409_),
    .X(_00410_));
 sky130_fd_sc_hd__clkbuf_1 _05127_ (.A(_00410_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _05128_ (.A0(_00293_),
    .A1(net4106),
    .S(_00409_),
    .X(_00411_));
 sky130_fd_sc_hd__clkbuf_1 _05129_ (.A(_00411_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _05130_ (.A0(_00295_),
    .A1(net3317),
    .S(_00409_),
    .X(_00412_));
 sky130_fd_sc_hd__clkbuf_1 _05131_ (.A(_00412_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _05132_ (.A0(_00297_),
    .A1(net3970),
    .S(_00409_),
    .X(_00413_));
 sky130_fd_sc_hd__clkbuf_1 _05133_ (.A(_00413_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[35] ));
 sky130_fd_sc_hd__clkbuf_4 _05134_ (.A(_00363_),
    .X(_00414_));
 sky130_fd_sc_hd__or2b_1 _05135_ (.A(_00327_),
    .B_N(_00313_),
    .X(_00415_));
 sky130_fd_sc_hd__or2_1 _05136_ (.A(_00325_),
    .B(_00406_),
    .X(_00416_));
 sky130_fd_sc_hd__nand2_1 _05137_ (.A(net4134),
    .B(_00416_),
    .Y(_00417_));
 sky130_fd_sc_hd__o31a_1 _05138_ (.A1(_00325_),
    .A2(_00329_),
    .A3(_00415_),
    .B1(_00417_),
    .X(_00418_));
 sky130_fd_sc_hd__o21ai_1 _05139_ (.A1(_00414_),
    .A2(_00418_),
    .B1(_00238_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[36] ));
 sky130_fd_sc_hd__nand2_1 _05140_ (.A(net3842),
    .B(_00416_),
    .Y(_00419_));
 sky130_fd_sc_hd__o31a_1 _05141_ (.A1(_00325_),
    .A2(_00335_),
    .A3(_00415_),
    .B1(_00419_),
    .X(_00420_));
 sky130_fd_sc_hd__o21ai_1 _05142_ (.A1(_00414_),
    .A2(_00420_),
    .B1(_00306_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[37] ));
 sky130_fd_sc_hd__nand2_1 _05143_ (.A(net4008),
    .B(_00416_),
    .Y(_00421_));
 sky130_fd_sc_hd__o31a_1 _05144_ (.A1(_00325_),
    .A2(_00338_),
    .A3(_00415_),
    .B1(_00421_),
    .X(_00422_));
 sky130_fd_sc_hd__o21ai_1 _05145_ (.A1(_00414_),
    .A2(_00422_),
    .B1(_00252_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[38] ));
 sky130_fd_sc_hd__nand2_1 _05146_ (.A(net3978),
    .B(_00416_),
    .Y(_00423_));
 sky130_fd_sc_hd__o31a_1 _05147_ (.A1(_00325_),
    .A2(_00341_),
    .A3(_00415_),
    .B1(_00423_),
    .X(_00424_));
 sky130_fd_sc_hd__clkbuf_8 _05148_ (.A(_00227_),
    .X(_00425_));
 sky130_fd_sc_hd__o21ai_1 _05149_ (.A1(_00414_),
    .A2(_00424_),
    .B1(_00425_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[39] ));
 sky130_fd_sc_hd__and3b_1 _05150_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[2].x.cfgd ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.cfgd ),
    .C(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ),
    .X(_00426_));
 sky130_fd_sc_hd__buf_2 _05151_ (.A(_00426_),
    .X(_00427_));
 sky130_fd_sc_hd__or2_1 _05152_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[3] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ),
    .X(_00428_));
 sky130_fd_sc_hd__or2_1 _05153_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ),
    .B(_00428_),
    .X(_00429_));
 sky130_fd_sc_hd__or2_1 _05154_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[5] ),
    .B(_00429_),
    .X(_00430_));
 sky130_fd_sc_hd__clkbuf_4 _05155_ (.A(_00430_),
    .X(_00431_));
 sky130_fd_sc_hd__inv_2 _05156_ (.A(_00431_),
    .Y(_00432_));
 sky130_fd_sc_hd__a21oi_4 _05157_ (.A1(_00427_),
    .A2(_00432_),
    .B1(_00267_),
    .Y(_00433_));
 sky130_fd_sc_hd__mux2_1 _05158_ (.A0(_00288_),
    .A1(net4123),
    .S(_00433_),
    .X(_00434_));
 sky130_fd_sc_hd__clkbuf_1 _05159_ (.A(_00434_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _05160_ (.A0(_00293_),
    .A1(net4098),
    .S(_00433_),
    .X(_00435_));
 sky130_fd_sc_hd__clkbuf_1 _05161_ (.A(_00435_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _05162_ (.A0(_00295_),
    .A1(net4188),
    .S(_00433_),
    .X(_00436_));
 sky130_fd_sc_hd__clkbuf_1 _05163_ (.A(_00436_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _05164_ (.A0(_00297_),
    .A1(net4211),
    .S(_00433_),
    .X(_00437_));
 sky130_fd_sc_hd__clkbuf_1 _05165_ (.A(_00437_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[3] ));
 sky130_fd_sc_hd__clkbuf_2 _05166_ (.A(net3749),
    .X(_00438_));
 sky130_fd_sc_hd__or3b_4 _05167_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ),
    .B(_00438_),
    .C_N(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ),
    .X(_00439_));
 sky130_fd_sc_hd__nand2_1 _05168_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[5] ),
    .B(_00429_),
    .Y(_00440_));
 sky130_fd_sc_hd__and2_1 _05169_ (.A(_00431_),
    .B(_00440_),
    .X(_00441_));
 sky130_fd_sc_hd__nand2_1 _05170_ (.A(_00427_),
    .B(_00441_),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_4 _05171_ (.A(_00170_),
    .B(_00431_),
    .Y(_00443_));
 sky130_fd_sc_hd__nor3b_1 _05172_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ),
    .B(_00438_),
    .C_N(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ),
    .Y(_00444_));
 sky130_fd_sc_hd__and3b_1 _05173_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[5] ),
    .B(_00427_),
    .C(_00444_),
    .X(_00445_));
 sky130_fd_sc_hd__inv_2 _05174_ (.A(net3743),
    .Y(_00446_));
 sky130_fd_sc_hd__o32a_1 _05175_ (.A1(_00439_),
    .A2(_00442_),
    .A3(_00443_),
    .B1(_00445_),
    .B2(_00446_),
    .X(_00447_));
 sky130_fd_sc_hd__buf_4 _05176_ (.A(_00237_),
    .X(_00448_));
 sky130_fd_sc_hd__o21ai_1 _05177_ (.A1(_00414_),
    .A2(_00447_),
    .B1(_00448_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[4] ));
 sky130_fd_sc_hd__nand2_4 _05178_ (.A(_00211_),
    .B(_00431_),
    .Y(_00449_));
 sky130_fd_sc_hd__inv_2 _05179_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ),
    .Y(_00450_));
 sky130_fd_sc_hd__o32a_1 _05180_ (.A1(_00439_),
    .A2(_00442_),
    .A3(_00449_),
    .B1(_00445_),
    .B2(_00450_),
    .X(_00451_));
 sky130_fd_sc_hd__o21ai_1 _05181_ (.A1(_00414_),
    .A2(_00451_),
    .B1(_00306_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[5] ));
 sky130_fd_sc_hd__nand2_2 _05182_ (.A(_00187_),
    .B(_00431_),
    .Y(_00452_));
 sky130_fd_sc_hd__inv_2 _05183_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ),
    .Y(_00453_));
 sky130_fd_sc_hd__o32a_1 _05184_ (.A1(_00439_),
    .A2(_00442_),
    .A3(_00452_),
    .B1(_00445_),
    .B2(_00453_),
    .X(_00454_));
 sky130_fd_sc_hd__o21ai_1 _05185_ (.A1(_00414_),
    .A2(_00454_),
    .B1(_00252_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[6] ));
 sky130_fd_sc_hd__nand2_4 _05186_ (.A(_00264_),
    .B(_00431_),
    .Y(_00455_));
 sky130_fd_sc_hd__inv_2 _05187_ (.A(net4083),
    .Y(_00456_));
 sky130_fd_sc_hd__o32a_1 _05188_ (.A1(_00439_),
    .A2(_00442_),
    .A3(_00455_),
    .B1(_00445_),
    .B2(_00456_),
    .X(_00457_));
 sky130_fd_sc_hd__o21ai_1 _05189_ (.A1(_00414_),
    .A2(_00457_),
    .B1(_00425_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _05190_ (.A(net3422),
    .Y(_00458_));
 sky130_fd_sc_hd__inv_2 _05191_ (.A(_00429_),
    .Y(_00459_));
 sky130_fd_sc_hd__and2_1 _05192_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ),
    .B(_00428_),
    .X(_00460_));
 sky130_fd_sc_hd__or4b_2 _05193_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[5] ),
    .B(_00459_),
    .C(_00460_),
    .D_N(_00426_),
    .X(_00461_));
 sky130_fd_sc_hd__or3b_2 _05194_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ),
    .B(_00461_),
    .C_N(_00438_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _05195_ (.A0(_00443_),
    .A1(_00458_),
    .S(_00462_),
    .X(_00463_));
 sky130_fd_sc_hd__o21ai_1 _05196_ (.A1(_00414_),
    .A2(_00463_),
    .B1(_00448_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[8] ));
 sky130_fd_sc_hd__inv_2 _05197_ (.A(net3941),
    .Y(_00464_));
 sky130_fd_sc_hd__mux2_1 _05198_ (.A0(_00449_),
    .A1(_00464_),
    .S(_00462_),
    .X(_00465_));
 sky130_fd_sc_hd__o21ai_1 _05199_ (.A1(_00414_),
    .A2(_00465_),
    .B1(_00306_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[9] ));
 sky130_fd_sc_hd__clkbuf_4 _05200_ (.A(_00363_),
    .X(_00466_));
 sky130_fd_sc_hd__inv_2 _05201_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ),
    .Y(_00467_));
 sky130_fd_sc_hd__mux2_1 _05202_ (.A0(_00452_),
    .A1(_00467_),
    .S(_00462_),
    .X(_00468_));
 sky130_fd_sc_hd__o21ai_1 _05203_ (.A1(_00466_),
    .A2(_00468_),
    .B1(_00252_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[10] ));
 sky130_fd_sc_hd__clkinv_2 _05204_ (.A(net4117),
    .Y(_00469_));
 sky130_fd_sc_hd__mux2_1 _05205_ (.A0(_00455_),
    .A1(_00469_),
    .S(_00462_),
    .X(_00470_));
 sky130_fd_sc_hd__o21ai_1 _05206_ (.A1(_00466_),
    .A2(_00470_),
    .B1(_00425_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[11] ));
 sky130_fd_sc_hd__inv_2 _05207_ (.A(net3926),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _05208_ (.A(_00438_),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ),
    .Y(_00472_));
 sky130_fd_sc_hd__nor2_2 _05209_ (.A(_00461_),
    .B(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__mux2_1 _05210_ (.A0(_00471_),
    .A1(_00443_),
    .S(_00473_),
    .X(_00474_));
 sky130_fd_sc_hd__o21ai_1 _05211_ (.A1(_00466_),
    .A2(_00474_),
    .B1(_00448_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[12] ));
 sky130_fd_sc_hd__inv_2 _05212_ (.A(net3683),
    .Y(_00475_));
 sky130_fd_sc_hd__mux2_1 _05213_ (.A0(_00475_),
    .A1(_00449_),
    .S(_00473_),
    .X(_00476_));
 sky130_fd_sc_hd__o21ai_1 _05214_ (.A1(_00466_),
    .A2(_00476_),
    .B1(_00306_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[13] ));
 sky130_fd_sc_hd__inv_2 _05215_ (.A(net3395),
    .Y(_00477_));
 sky130_fd_sc_hd__mux2_1 _05216_ (.A0(_00477_),
    .A1(_00452_),
    .S(_00473_),
    .X(_00478_));
 sky130_fd_sc_hd__buf_4 _05217_ (.A(_00251_),
    .X(_00479_));
 sky130_fd_sc_hd__o21ai_1 _05218_ (.A1(_00466_),
    .A2(_00478_),
    .B1(_00479_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[14] ));
 sky130_fd_sc_hd__inv_2 _05219_ (.A(net4054),
    .Y(_00480_));
 sky130_fd_sc_hd__mux2_1 _05220_ (.A0(_00480_),
    .A1(_00455_),
    .S(_00473_),
    .X(_00481_));
 sky130_fd_sc_hd__o21ai_1 _05221_ (.A1(_00466_),
    .A2(_00481_),
    .B1(_00425_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[15] ));
 sky130_fd_sc_hd__nor2_4 _05222_ (.A(_00428_),
    .B(_00461_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _05223_ (.A(_00443_),
    .B(_00482_),
    .Y(_00483_));
 sky130_fd_sc_hd__or2_1 _05224_ (.A(net4193),
    .B(_00482_),
    .X(_00484_));
 sky130_fd_sc_hd__a31o_1 _05225_ (.A1(_00367_),
    .A2(_00483_),
    .A3(_00484_),
    .B1(_00210_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _05226_ (.A(_00449_),
    .B(_00482_),
    .Y(_00485_));
 sky130_fd_sc_hd__or2_1 _05227_ (.A(net4133),
    .B(_00482_),
    .X(_00486_));
 sky130_fd_sc_hd__buf_6 _05228_ (.A(_00215_),
    .X(_00487_));
 sky130_fd_sc_hd__a31o_1 _05229_ (.A1(_00367_),
    .A2(_00485_),
    .A3(_00486_),
    .B1(_00487_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _05230_ (.A(_00452_),
    .B(_00482_),
    .Y(_00488_));
 sky130_fd_sc_hd__or2_1 _05231_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[18] ),
    .B(_00482_),
    .X(_00489_));
 sky130_fd_sc_hd__a31o_1 _05232_ (.A1(_00367_),
    .A2(_00488_),
    .A3(_00489_),
    .B1(_00394_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _05233_ (.A(net3433),
    .B(_00482_),
    .Y(_00490_));
 sky130_fd_sc_hd__a211o_1 _05234_ (.A1(_00455_),
    .A2(_00482_),
    .B1(_00490_),
    .C1(_00268_),
    .X(_00491_));
 sky130_fd_sc_hd__nand2_1 _05235_ (.A(_00263_),
    .B(_00491_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[19] ));
 sky130_fd_sc_hd__inv_2 _05236_ (.A(net4120),
    .Y(_00492_));
 sky130_fd_sc_hd__and3_1 _05237_ (.A(_00427_),
    .B(_00431_),
    .C(_00440_),
    .X(_00493_));
 sky130_fd_sc_hd__and4b_2 _05238_ (.A_N(_00438_),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ),
    .C(_00493_),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _05239_ (.A0(_00492_),
    .A1(_00443_),
    .S(_00494_),
    .X(_00495_));
 sky130_fd_sc_hd__o21ai_1 _05240_ (.A1(_00466_),
    .A2(_00495_),
    .B1(_00448_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[20] ));
 sky130_fd_sc_hd__or2_1 _05241_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[21] ),
    .B(_00494_),
    .X(_00496_));
 sky130_fd_sc_hd__nand2_1 _05242_ (.A(_00449_),
    .B(_00494_),
    .Y(_00497_));
 sky130_fd_sc_hd__a31o_1 _05243_ (.A1(_00367_),
    .A2(_00496_),
    .A3(_00497_),
    .B1(_00487_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[21] ));
 sky130_fd_sc_hd__inv_2 _05244_ (.A(net4028),
    .Y(_00498_));
 sky130_fd_sc_hd__mux2_1 _05245_ (.A0(_00498_),
    .A1(_00452_),
    .S(_00494_),
    .X(_00499_));
 sky130_fd_sc_hd__o21ai_1 _05246_ (.A1(_00466_),
    .A2(_00499_),
    .B1(_00479_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[22] ));
 sky130_fd_sc_hd__inv_2 _05247_ (.A(net3984),
    .Y(_00500_));
 sky130_fd_sc_hd__mux2_1 _05248_ (.A0(_00500_),
    .A1(_00455_),
    .S(_00494_),
    .X(_00501_));
 sky130_fd_sc_hd__o21ai_1 _05249_ (.A1(_00466_),
    .A2(_00501_),
    .B1(_00425_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[23] ));
 sky130_fd_sc_hd__inv_2 _05250_ (.A(net3256),
    .Y(_00502_));
 sky130_fd_sc_hd__and4b_2 _05251_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ),
    .B(_00493_),
    .C(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ),
    .D(_00438_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _05252_ (.A0(_00502_),
    .A1(_00443_),
    .S(_00503_),
    .X(_00504_));
 sky130_fd_sc_hd__o21ai_1 _05253_ (.A1(_00466_),
    .A2(_00504_),
    .B1(_00448_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[24] ));
 sky130_fd_sc_hd__clkbuf_4 _05254_ (.A(_00363_),
    .X(_00505_));
 sky130_fd_sc_hd__inv_2 _05255_ (.A(net4070),
    .Y(_00506_));
 sky130_fd_sc_hd__mux2_1 _05256_ (.A0(_00506_),
    .A1(_00449_),
    .S(_00503_),
    .X(_00507_));
 sky130_fd_sc_hd__buf_4 _05257_ (.A(_00305_),
    .X(_00508_));
 sky130_fd_sc_hd__o21ai_1 _05258_ (.A1(_00505_),
    .A2(_00507_),
    .B1(_00508_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[25] ));
 sky130_fd_sc_hd__nand2_1 _05259_ (.A(_00452_),
    .B(_00503_),
    .Y(_00509_));
 sky130_fd_sc_hd__or2_1 _05260_ (.A(net4166),
    .B(_00503_),
    .X(_00510_));
 sky130_fd_sc_hd__a31o_1 _05261_ (.A1(_00367_),
    .A2(_00509_),
    .A3(_00510_),
    .B1(_00394_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[26] ));
 sky130_fd_sc_hd__inv_2 _05262_ (.A(net3925),
    .Y(_00511_));
 sky130_fd_sc_hd__mux2_1 _05263_ (.A0(_00511_),
    .A1(_00455_),
    .S(_00503_),
    .X(_00512_));
 sky130_fd_sc_hd__o21ai_1 _05264_ (.A1(_00505_),
    .A2(_00512_),
    .B1(_00425_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[27] ));
 sky130_fd_sc_hd__inv_2 _05265_ (.A(net4027),
    .Y(_00513_));
 sky130_fd_sc_hd__and4_2 _05266_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ),
    .B(_00438_),
    .C(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ),
    .D(_00493_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _05267_ (.A0(_00513_),
    .A1(_00443_),
    .S(_00514_),
    .X(_00515_));
 sky130_fd_sc_hd__o21ai_1 _05268_ (.A1(_00505_),
    .A2(_00515_),
    .B1(_00448_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[28] ));
 sky130_fd_sc_hd__inv_2 _05269_ (.A(net3309),
    .Y(_00516_));
 sky130_fd_sc_hd__mux2_1 _05270_ (.A0(_00516_),
    .A1(_00449_),
    .S(_00514_),
    .X(_00517_));
 sky130_fd_sc_hd__o21ai_1 _05271_ (.A1(_00505_),
    .A2(_00517_),
    .B1(_00508_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[29] ));
 sky130_fd_sc_hd__inv_2 _05272_ (.A(net3650),
    .Y(_00518_));
 sky130_fd_sc_hd__mux2_1 _05273_ (.A0(_00518_),
    .A1(_00452_),
    .S(_00514_),
    .X(_00519_));
 sky130_fd_sc_hd__o21ai_1 _05274_ (.A1(_00505_),
    .A2(_00519_),
    .B1(_00479_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[30] ));
 sky130_fd_sc_hd__nor2_1 _05275_ (.A(net3968),
    .B(_00514_),
    .Y(_00520_));
 sky130_fd_sc_hd__a211o_1 _05276_ (.A1(_00455_),
    .A2(_00514_),
    .B1(_00520_),
    .C1(_00268_),
    .X(_00521_));
 sky130_fd_sc_hd__nand2_1 _05277_ (.A(_00263_),
    .B(_00521_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[31] ));
 sky130_fd_sc_hd__buf_6 _05278_ (.A(_00180_),
    .X(_00522_));
 sky130_fd_sc_hd__a31o_2 _05279_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[5] ),
    .A2(_00427_),
    .A3(_00459_),
    .B1(_00522_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _05280_ (.A0(net4096),
    .A1(_00172_),
    .S(_00523_),
    .X(_00524_));
 sky130_fd_sc_hd__clkbuf_1 _05281_ (.A(_00524_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _05282_ (.A0(net4102),
    .A1(_00185_),
    .S(_00523_),
    .X(_00525_));
 sky130_fd_sc_hd__clkbuf_1 _05283_ (.A(_00525_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _05284_ (.A0(net4214),
    .A1(_00189_),
    .S(_00523_),
    .X(_00526_));
 sky130_fd_sc_hd__clkbuf_1 _05285_ (.A(_00526_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[34] ));
 sky130_fd_sc_hd__buf_6 _05286_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ),
    .X(_00527_));
 sky130_fd_sc_hd__buf_8 _05287_ (.A(_00527_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _05288_ (.A0(net4203),
    .A1(_00528_),
    .S(_00523_),
    .X(_00529_));
 sky130_fd_sc_hd__clkbuf_1 _05289_ (.A(_00529_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2b_1 _05290_ (.A(_00441_),
    .B_N(_00427_),
    .X(_00530_));
 sky130_fd_sc_hd__and3_1 _05291_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[5] ),
    .B(_00427_),
    .C(_00444_),
    .X(_00531_));
 sky130_fd_sc_hd__inv_2 _05292_ (.A(net4113),
    .Y(_00532_));
 sky130_fd_sc_hd__o32a_1 _05293_ (.A1(_00439_),
    .A2(_00443_),
    .A3(_00530_),
    .B1(_00531_),
    .B2(_00532_),
    .X(_00533_));
 sky130_fd_sc_hd__o21ai_1 _05294_ (.A1(_00505_),
    .A2(_00533_),
    .B1(_00448_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[36] ));
 sky130_fd_sc_hd__inv_2 _05295_ (.A(net3538),
    .Y(_00534_));
 sky130_fd_sc_hd__o32a_1 _05296_ (.A1(_00439_),
    .A2(_00449_),
    .A3(_00530_),
    .B1(_00531_),
    .B2(_00534_),
    .X(_00535_));
 sky130_fd_sc_hd__o21ai_1 _05297_ (.A1(_00505_),
    .A2(_00535_),
    .B1(_00508_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[37] ));
 sky130_fd_sc_hd__inv_2 _05298_ (.A(net3811),
    .Y(_00536_));
 sky130_fd_sc_hd__o32a_1 _05299_ (.A1(_00439_),
    .A2(_00452_),
    .A3(_00530_),
    .B1(_00531_),
    .B2(_00536_),
    .X(_00537_));
 sky130_fd_sc_hd__o21ai_1 _05300_ (.A1(_00505_),
    .A2(_00537_),
    .B1(_00479_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[38] ));
 sky130_fd_sc_hd__inv_2 _05301_ (.A(net3504),
    .Y(_00538_));
 sky130_fd_sc_hd__o32a_1 _05302_ (.A1(_00439_),
    .A2(_00455_),
    .A3(_00530_),
    .B1(_00531_),
    .B2(_00538_),
    .X(_00539_));
 sky130_fd_sc_hd__o21ai_1 _05303_ (.A1(_00505_),
    .A2(_00539_),
    .B1(_00425_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[39] ));
 sky130_fd_sc_hd__buf_4 _05304_ (.A(_00171_),
    .X(_00540_));
 sky130_fd_sc_hd__and3b_1 _05305_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[3].x.cfgd ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.cfgd ),
    .C(_00311_),
    .X(_00541_));
 sky130_fd_sc_hd__buf_2 _05306_ (.A(_00541_),
    .X(_00542_));
 sky130_fd_sc_hd__or3_1 _05307_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[3] ),
    .C(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[2] ),
    .X(_00543_));
 sky130_fd_sc_hd__or2_1 _05308_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[5] ),
    .B(_00543_),
    .X(_00544_));
 sky130_fd_sc_hd__clkbuf_4 _05309_ (.A(_00544_),
    .X(_00545_));
 sky130_fd_sc_hd__inv_2 _05310_ (.A(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__a21oi_2 _05311_ (.A1(_00542_),
    .A2(_00546_),
    .B1(_00267_),
    .Y(_00547_));
 sky130_fd_sc_hd__mux2_1 _05312_ (.A0(_00540_),
    .A1(net4163),
    .S(_00547_),
    .X(_00548_));
 sky130_fd_sc_hd__clkbuf_1 _05313_ (.A(_00548_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[0] ));
 sky130_fd_sc_hd__buf_4 _05314_ (.A(_00184_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _05315_ (.A0(_00549_),
    .A1(net4207),
    .S(_00547_),
    .X(_00550_));
 sky130_fd_sc_hd__clkbuf_1 _05316_ (.A(_00550_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[1] ));
 sky130_fd_sc_hd__buf_8 _05317_ (.A(_00187_),
    .X(_00551_));
 sky130_fd_sc_hd__buf_4 _05318_ (.A(_00551_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _05319_ (.A0(_00552_),
    .A1(net3914),
    .S(_00547_),
    .X(_00553_));
 sky130_fd_sc_hd__clkbuf_1 _05320_ (.A(_00553_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _05321_ (.A0(_00297_),
    .A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ),
    .S(_00547_),
    .X(_00554_));
 sky130_fd_sc_hd__clkbuf_1 _05322_ (.A(_00554_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[3] ));
 sky130_fd_sc_hd__clkbuf_2 _05323_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[3] ),
    .X(_00555_));
 sky130_fd_sc_hd__clkbuf_2 _05324_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[2] ),
    .X(_00556_));
 sky130_fd_sc_hd__or3b_1 _05325_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ),
    .B(_00555_),
    .C_N(_00556_),
    .X(_00557_));
 sky130_fd_sc_hd__buf_2 _05326_ (.A(_00557_),
    .X(_00558_));
 sky130_fd_sc_hd__nand2_1 _05327_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[5] ),
    .B(_00543_),
    .Y(_00559_));
 sky130_fd_sc_hd__and2_1 _05328_ (.A(_00545_),
    .B(_00559_),
    .X(_00560_));
 sky130_fd_sc_hd__nand2_1 _05329_ (.A(_00542_),
    .B(_00560_),
    .Y(_00561_));
 sky130_fd_sc_hd__nand2_2 _05330_ (.A(_00170_),
    .B(_00545_),
    .Y(_00562_));
 sky130_fd_sc_hd__nor3b_1 _05331_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[3] ),
    .C_N(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[2] ),
    .Y(_00563_));
 sky130_fd_sc_hd__and3b_1 _05332_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[5] ),
    .B(_00542_),
    .C(_00563_),
    .X(_00564_));
 sky130_fd_sc_hd__inv_2 _05333_ (.A(net3688),
    .Y(_00565_));
 sky130_fd_sc_hd__o32a_1 _05334_ (.A1(_00558_),
    .A2(_00561_),
    .A3(_00562_),
    .B1(_00564_),
    .B2(_00565_),
    .X(_00566_));
 sky130_fd_sc_hd__o21ai_1 _05335_ (.A1(_00505_),
    .A2(_00566_),
    .B1(_00448_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[4] ));
 sky130_fd_sc_hd__buf_2 _05336_ (.A(_00363_),
    .X(_00567_));
 sky130_fd_sc_hd__nand2_4 _05337_ (.A(_00211_),
    .B(_00545_),
    .Y(_00568_));
 sky130_fd_sc_hd__inv_2 _05338_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ),
    .Y(_00569_));
 sky130_fd_sc_hd__o32a_1 _05339_ (.A1(_00558_),
    .A2(_00561_),
    .A3(_00568_),
    .B1(_00564_),
    .B2(_00569_),
    .X(_00570_));
 sky130_fd_sc_hd__o21ai_1 _05340_ (.A1(_00567_),
    .A2(_00570_),
    .B1(_00508_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[5] ));
 sky130_fd_sc_hd__nand2_4 _05341_ (.A(_00187_),
    .B(_00545_),
    .Y(_00571_));
 sky130_fd_sc_hd__inv_2 _05342_ (.A(net4107),
    .Y(_00572_));
 sky130_fd_sc_hd__o32a_1 _05343_ (.A1(_00558_),
    .A2(_00561_),
    .A3(_00571_),
    .B1(_00564_),
    .B2(_00572_),
    .X(_00573_));
 sky130_fd_sc_hd__o21ai_1 _05344_ (.A1(_00567_),
    .A2(_00573_),
    .B1(_00479_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[6] ));
 sky130_fd_sc_hd__nand2_4 _05345_ (.A(_00264_),
    .B(_00545_),
    .Y(_00574_));
 sky130_fd_sc_hd__inv_2 _05346_ (.A(net4068),
    .Y(_00575_));
 sky130_fd_sc_hd__o32a_1 _05347_ (.A1(_00558_),
    .A2(_00561_),
    .A3(_00574_),
    .B1(_00564_),
    .B2(_00575_),
    .X(_00576_));
 sky130_fd_sc_hd__o21ai_1 _05348_ (.A1(_00567_),
    .A2(_00576_),
    .B1(_00425_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _05349_ (.A(net4037),
    .Y(_00577_));
 sky130_fd_sc_hd__o21a_1 _05350_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[3] ),
    .A2(_00556_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ),
    .X(_00578_));
 sky130_fd_sc_hd__or4bb_2 _05351_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[5] ),
    .B(_00578_),
    .C_N(_00541_),
    .D_N(_00543_),
    .X(_00579_));
 sky130_fd_sc_hd__or3b_2 _05352_ (.A(_00556_),
    .B(_00579_),
    .C_N(_00555_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _05353_ (.A0(_00562_),
    .A1(_00577_),
    .S(_00580_),
    .X(_00581_));
 sky130_fd_sc_hd__o21ai_1 _05354_ (.A1(_00567_),
    .A2(_00581_),
    .B1(_00448_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[8] ));
 sky130_fd_sc_hd__inv_2 _05355_ (.A(net3287),
    .Y(_00582_));
 sky130_fd_sc_hd__mux2_1 _05356_ (.A0(_00568_),
    .A1(_00582_),
    .S(_00580_),
    .X(_00583_));
 sky130_fd_sc_hd__o21ai_1 _05357_ (.A1(_00567_),
    .A2(_00583_),
    .B1(_00508_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[9] ));
 sky130_fd_sc_hd__inv_2 _05358_ (.A(net4145),
    .Y(_00584_));
 sky130_fd_sc_hd__mux2_1 _05359_ (.A0(_00571_),
    .A1(_00584_),
    .S(_00580_),
    .X(_00585_));
 sky130_fd_sc_hd__o21ai_1 _05360_ (.A1(_00567_),
    .A2(_00585_),
    .B1(_00479_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[10] ));
 sky130_fd_sc_hd__clkinv_2 _05361_ (.A(net4015),
    .Y(_00586_));
 sky130_fd_sc_hd__mux2_1 _05362_ (.A0(_00574_),
    .A1(_00586_),
    .S(_00580_),
    .X(_00587_));
 sky130_fd_sc_hd__o21ai_1 _05363_ (.A1(_00567_),
    .A2(_00587_),
    .B1(_00425_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[11] ));
 sky130_fd_sc_hd__inv_2 _05364_ (.A(net3882),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _05365_ (.A(_00555_),
    .B(_00556_),
    .Y(_00589_));
 sky130_fd_sc_hd__nor2_2 _05366_ (.A(_00579_),
    .B(_00589_),
    .Y(_00590_));
 sky130_fd_sc_hd__mux2_1 _05367_ (.A0(_00588_),
    .A1(_00562_),
    .S(_00590_),
    .X(_00591_));
 sky130_fd_sc_hd__o21ai_1 _05368_ (.A1(_00567_),
    .A2(_00591_),
    .B1(_00448_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[12] ));
 sky130_fd_sc_hd__inv_2 _05369_ (.A(net3946),
    .Y(_00592_));
 sky130_fd_sc_hd__mux2_1 _05370_ (.A0(_00592_),
    .A1(_00568_),
    .S(_00590_),
    .X(_00593_));
 sky130_fd_sc_hd__o21ai_1 _05371_ (.A1(_00567_),
    .A2(_00593_),
    .B1(_00508_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[13] ));
 sky130_fd_sc_hd__inv_2 _05372_ (.A(net3474),
    .Y(_00594_));
 sky130_fd_sc_hd__mux2_1 _05373_ (.A0(_00594_),
    .A1(_00571_),
    .S(_00590_),
    .X(_00595_));
 sky130_fd_sc_hd__o21ai_1 _05374_ (.A1(_00567_),
    .A2(_00595_),
    .B1(_00479_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[14] ));
 sky130_fd_sc_hd__clkbuf_4 _05375_ (.A(_00363_),
    .X(_00596_));
 sky130_fd_sc_hd__inv_2 _05376_ (.A(net3185),
    .Y(_00597_));
 sky130_fd_sc_hd__mux2_1 _05377_ (.A0(_00597_),
    .A1(_00574_),
    .S(_00590_),
    .X(_00598_));
 sky130_fd_sc_hd__o21ai_1 _05378_ (.A1(_00596_),
    .A2(_00598_),
    .B1(_00425_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[15] ));
 sky130_fd_sc_hd__clkbuf_4 _05379_ (.A(_00196_),
    .X(_00599_));
 sky130_fd_sc_hd__nor3_2 _05380_ (.A(_00555_),
    .B(_00556_),
    .C(_00579_),
    .Y(_00600_));
 sky130_fd_sc_hd__nand2_1 _05381_ (.A(_00562_),
    .B(_00600_),
    .Y(_00601_));
 sky130_fd_sc_hd__or2_1 _05382_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ),
    .B(_00600_),
    .X(_00602_));
 sky130_fd_sc_hd__buf_6 _05383_ (.A(_00208_),
    .X(_00603_));
 sky130_fd_sc_hd__a31o_1 _05384_ (.A1(_00599_),
    .A2(_00601_),
    .A3(_00602_),
    .B1(_00603_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _05385_ (.A(_00568_),
    .B(_00600_),
    .Y(_00604_));
 sky130_fd_sc_hd__or2_1 _05386_ (.A(net4104),
    .B(_00600_),
    .X(_00605_));
 sky130_fd_sc_hd__a31o_1 _05387_ (.A1(_00599_),
    .A2(_00604_),
    .A3(_00605_),
    .B1(_00487_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _05388_ (.A(_00571_),
    .B(_00600_),
    .Y(_00606_));
 sky130_fd_sc_hd__or2_1 _05389_ (.A(net4064),
    .B(_00600_),
    .X(_00607_));
 sky130_fd_sc_hd__a31o_1 _05390_ (.A1(_00599_),
    .A2(_00606_),
    .A3(_00607_),
    .B1(_00394_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _05391_ (.A(net3890),
    .B(_00600_),
    .Y(_00608_));
 sky130_fd_sc_hd__a211o_1 _05392_ (.A1(_00574_),
    .A2(_00600_),
    .B1(_00608_),
    .C1(_00268_),
    .X(_00609_));
 sky130_fd_sc_hd__nand2_1 _05393_ (.A(_00263_),
    .B(_00609_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[19] ));
 sky130_fd_sc_hd__inv_2 _05394_ (.A(net4196),
    .Y(_00610_));
 sky130_fd_sc_hd__and3_1 _05395_ (.A(_00542_),
    .B(_00545_),
    .C(_00559_),
    .X(_00611_));
 sky130_fd_sc_hd__and4b_2 _05396_ (.A_N(_00555_),
    .B(_00556_),
    .C(_00611_),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _05397_ (.A0(_00610_),
    .A1(_00562_),
    .S(_00612_),
    .X(_00613_));
 sky130_fd_sc_hd__buf_4 _05398_ (.A(_00237_),
    .X(_00614_));
 sky130_fd_sc_hd__o21ai_1 _05399_ (.A1(_00596_),
    .A2(_00613_),
    .B1(_00614_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[20] ));
 sky130_fd_sc_hd__or2_1 _05400_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ),
    .B(_00612_),
    .X(_00615_));
 sky130_fd_sc_hd__nand2_1 _05401_ (.A(_00568_),
    .B(_00612_),
    .Y(_00616_));
 sky130_fd_sc_hd__a31o_1 _05402_ (.A1(_00599_),
    .A2(_00615_),
    .A3(_00616_),
    .B1(_00487_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[21] ));
 sky130_fd_sc_hd__inv_2 _05403_ (.A(net3282),
    .Y(_00617_));
 sky130_fd_sc_hd__mux2_1 _05404_ (.A0(_00617_),
    .A1(_00571_),
    .S(_00612_),
    .X(_00618_));
 sky130_fd_sc_hd__o21ai_1 _05405_ (.A1(_00596_),
    .A2(_00618_),
    .B1(_00479_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[22] ));
 sky130_fd_sc_hd__inv_2 _05406_ (.A(net4006),
    .Y(_00619_));
 sky130_fd_sc_hd__mux2_1 _05407_ (.A0(_00619_),
    .A1(_00574_),
    .S(_00612_),
    .X(_00620_));
 sky130_fd_sc_hd__clkbuf_8 _05408_ (.A(_00226_),
    .X(_00621_));
 sky130_fd_sc_hd__o21ai_1 _05409_ (.A1(_00596_),
    .A2(_00620_),
    .B1(_00621_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[23] ));
 sky130_fd_sc_hd__inv_2 _05410_ (.A(net3715),
    .Y(_00622_));
 sky130_fd_sc_hd__and4b_2 _05411_ (.A_N(_00556_),
    .B(_00611_),
    .C(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ),
    .D(_00555_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _05412_ (.A0(_00622_),
    .A1(_00562_),
    .S(_00623_),
    .X(_00624_));
 sky130_fd_sc_hd__o21ai_1 _05413_ (.A1(_00596_),
    .A2(_00624_),
    .B1(_00614_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[24] ));
 sky130_fd_sc_hd__inv_2 _05414_ (.A(net4103),
    .Y(_00625_));
 sky130_fd_sc_hd__mux2_1 _05415_ (.A0(_00625_),
    .A1(_00568_),
    .S(_00623_),
    .X(_00626_));
 sky130_fd_sc_hd__o21ai_1 _05416_ (.A1(_00596_),
    .A2(_00626_),
    .B1(_00508_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[25] ));
 sky130_fd_sc_hd__or2_1 _05417_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ),
    .B(_00623_),
    .X(_00627_));
 sky130_fd_sc_hd__nand2_1 _05418_ (.A(_00571_),
    .B(_00623_),
    .Y(_00628_));
 sky130_fd_sc_hd__a31o_1 _05419_ (.A1(_00599_),
    .A2(_00627_),
    .A3(_00628_),
    .B1(_00394_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[26] ));
 sky130_fd_sc_hd__inv_2 _05420_ (.A(net3994),
    .Y(_00629_));
 sky130_fd_sc_hd__mux2_1 _05421_ (.A0(_00629_),
    .A1(_00574_),
    .S(_00623_),
    .X(_00630_));
 sky130_fd_sc_hd__o21ai_1 _05422_ (.A1(_00596_),
    .A2(_00630_),
    .B1(_00621_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[27] ));
 sky130_fd_sc_hd__inv_2 _05423_ (.A(net3738),
    .Y(_00631_));
 sky130_fd_sc_hd__and4_2 _05424_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ),
    .B(_00555_),
    .C(_00556_),
    .D(_00611_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _05425_ (.A0(_00631_),
    .A1(_00562_),
    .S(_00632_),
    .X(_00633_));
 sky130_fd_sc_hd__o21ai_1 _05426_ (.A1(_00596_),
    .A2(_00633_),
    .B1(_00614_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[28] ));
 sky130_fd_sc_hd__inv_2 _05427_ (.A(net3598),
    .Y(_00634_));
 sky130_fd_sc_hd__mux2_1 _05428_ (.A0(_00634_),
    .A1(_00568_),
    .S(_00632_),
    .X(_00635_));
 sky130_fd_sc_hd__o21ai_1 _05429_ (.A1(_00596_),
    .A2(_00635_),
    .B1(_00508_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[29] ));
 sky130_fd_sc_hd__inv_2 _05430_ (.A(net4043),
    .Y(_00636_));
 sky130_fd_sc_hd__mux2_1 _05431_ (.A0(_00636_),
    .A1(_00571_),
    .S(_00632_),
    .X(_00637_));
 sky130_fd_sc_hd__o21ai_1 _05432_ (.A1(_00596_),
    .A2(_00637_),
    .B1(_00479_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[30] ));
 sky130_fd_sc_hd__nor2_1 _05433_ (.A(net4086),
    .B(_00632_),
    .Y(_00638_));
 sky130_fd_sc_hd__a211o_1 _05434_ (.A1(_00574_),
    .A2(_00632_),
    .B1(_00638_),
    .C1(_00268_),
    .X(_00639_));
 sky130_fd_sc_hd__nand2_1 _05435_ (.A(_00263_),
    .B(_00639_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[31] ));
 sky130_fd_sc_hd__nand2_1 _05436_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[5] ),
    .B(_00542_),
    .Y(_00640_));
 sky130_fd_sc_hd__o21a_1 _05437_ (.A1(_00543_),
    .A2(_00640_),
    .B1(_00408_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _05438_ (.A0(_00540_),
    .A1(net4057),
    .S(_00641_),
    .X(_00642_));
 sky130_fd_sc_hd__clkbuf_1 _05439_ (.A(_00642_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _05440_ (.A0(_00549_),
    .A1(net3826),
    .S(_00641_),
    .X(_00643_));
 sky130_fd_sc_hd__clkbuf_1 _05441_ (.A(_00643_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _05442_ (.A0(_00552_),
    .A1(net3724),
    .S(_00641_),
    .X(_00644_));
 sky130_fd_sc_hd__clkbuf_1 _05443_ (.A(_00644_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _05444_ (.A0(_00297_),
    .A1(net4062),
    .S(_00641_),
    .X(_00645_));
 sky130_fd_sc_hd__clkbuf_1 _05445_ (.A(_00645_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[35] ));
 sky130_fd_sc_hd__clkbuf_4 _05446_ (.A(_00363_),
    .X(_00646_));
 sky130_fd_sc_hd__or2b_1 _05447_ (.A(_00560_),
    .B_N(_00542_),
    .X(_00647_));
 sky130_fd_sc_hd__nor2_1 _05448_ (.A(_00558_),
    .B(_00640_),
    .Y(_00648_));
 sky130_fd_sc_hd__inv_2 _05449_ (.A(net4205),
    .Y(_00649_));
 sky130_fd_sc_hd__o32a_1 _05450_ (.A1(_00558_),
    .A2(_00562_),
    .A3(_00647_),
    .B1(_00648_),
    .B2(_00649_),
    .X(_00650_));
 sky130_fd_sc_hd__o21ai_1 _05451_ (.A1(_00646_),
    .A2(_00650_),
    .B1(_00614_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[36] ));
 sky130_fd_sc_hd__inv_2 _05452_ (.A(net4069),
    .Y(_00651_));
 sky130_fd_sc_hd__o32a_1 _05453_ (.A1(_00558_),
    .A2(_00568_),
    .A3(_00647_),
    .B1(_00648_),
    .B2(_00651_),
    .X(_00652_));
 sky130_fd_sc_hd__o21ai_1 _05454_ (.A1(_00646_),
    .A2(_00652_),
    .B1(_00508_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[37] ));
 sky130_fd_sc_hd__inv_2 _05455_ (.A(net4095),
    .Y(_00653_));
 sky130_fd_sc_hd__o32a_1 _05456_ (.A1(_00558_),
    .A2(_00571_),
    .A3(_00647_),
    .B1(_00648_),
    .B2(_00653_),
    .X(_00654_));
 sky130_fd_sc_hd__o21ai_1 _05457_ (.A1(_00646_),
    .A2(_00654_),
    .B1(_00479_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[38] ));
 sky130_fd_sc_hd__inv_2 _05458_ (.A(net3307),
    .Y(_00655_));
 sky130_fd_sc_hd__o32a_1 _05459_ (.A1(_00558_),
    .A2(_00574_),
    .A3(_00647_),
    .B1(_00648_),
    .B2(_00655_),
    .X(_00656_));
 sky130_fd_sc_hd__o21ai_1 _05460_ (.A1(_00646_),
    .A2(_00656_),
    .B1(_00621_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[39] ));
 sky130_fd_sc_hd__clkinv_2 _05461_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ),
    .Y(_00657_));
 sky130_fd_sc_hd__clkinv_2 _05462_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[2] ),
    .Y(_00658_));
 sky130_fd_sc_hd__and3b_1 _05463_ (.A_N(net27),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.cfgd ),
    .C(_00311_),
    .X(_00659_));
 sky130_fd_sc_hd__clkbuf_4 _05464_ (.A(_00659_),
    .X(_00660_));
 sky130_fd_sc_hd__and2b_1 _05465_ (.A_N(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[4] ),
    .B(_00660_),
    .X(_00661_));
 sky130_fd_sc_hd__a31oi_4 _05466_ (.A1(_00657_),
    .A2(_00658_),
    .A3(_00661_),
    .B1(_00181_),
    .Y(_00662_));
 sky130_fd_sc_hd__mux2_1 _05467_ (.A0(_00540_),
    .A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[0] ),
    .S(_00662_),
    .X(_00663_));
 sky130_fd_sc_hd__clkbuf_1 _05468_ (.A(_00663_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _05469_ (.A0(_00549_),
    .A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[1] ),
    .S(_00662_),
    .X(_00664_));
 sky130_fd_sc_hd__clkbuf_1 _05470_ (.A(_00664_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _05471_ (.A0(_00552_),
    .A1(net3923),
    .S(_00662_),
    .X(_00665_));
 sky130_fd_sc_hd__clkbuf_1 _05472_ (.A(_00665_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _05473_ (.A0(_00297_),
    .A1(net3225),
    .S(_00662_),
    .X(_00666_));
 sky130_fd_sc_hd__clkbuf_1 _05474_ (.A(_00666_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[3] ));
 sky130_fd_sc_hd__a31o_2 _05475_ (.A1(_00657_),
    .A2(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[2] ),
    .A3(_00661_),
    .B1(_00522_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _05476_ (.A0(net4184),
    .A1(_00172_),
    .S(_00667_),
    .X(_00668_));
 sky130_fd_sc_hd__clkbuf_1 _05477_ (.A(_00668_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _05478_ (.A0(net4010),
    .A1(_00185_),
    .S(_00667_),
    .X(_00669_));
 sky130_fd_sc_hd__clkbuf_1 _05479_ (.A(_00669_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _05480_ (.A0(net3774),
    .A1(_00189_),
    .S(_00667_),
    .X(_00670_));
 sky130_fd_sc_hd__clkbuf_1 _05481_ (.A(_00670_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _05482_ (.A0(net3215),
    .A1(_00528_),
    .S(_00667_),
    .X(_00671_));
 sky130_fd_sc_hd__clkbuf_1 _05483_ (.A(_00671_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[7] ));
 sky130_fd_sc_hd__a31o_2 _05484_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ),
    .A2(_00658_),
    .A3(_00661_),
    .B1(_00522_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _05485_ (.A0(net4112),
    .A1(_00172_),
    .S(_00672_),
    .X(_00673_));
 sky130_fd_sc_hd__clkbuf_1 _05486_ (.A(_00673_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[8] ));
 sky130_fd_sc_hd__mux2_1 _05487_ (.A0(net3916),
    .A1(_00185_),
    .S(_00672_),
    .X(_00674_));
 sky130_fd_sc_hd__clkbuf_1 _05488_ (.A(_00674_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[9] ));
 sky130_fd_sc_hd__mux2_1 _05489_ (.A0(net3933),
    .A1(_00189_),
    .S(_00672_),
    .X(_00675_));
 sky130_fd_sc_hd__clkbuf_1 _05490_ (.A(_00675_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[10] ));
 sky130_fd_sc_hd__mux2_1 _05491_ (.A0(net3388),
    .A1(_00528_),
    .S(_00672_),
    .X(_00676_));
 sky130_fd_sc_hd__clkbuf_1 _05492_ (.A(_00676_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[11] ));
 sky130_fd_sc_hd__a31o_2 _05493_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ),
    .A2(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[2] ),
    .A3(_00661_),
    .B1(_00522_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _05494_ (.A0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ),
    .A1(_00172_),
    .S(_00677_),
    .X(_00678_));
 sky130_fd_sc_hd__clkbuf_1 _05495_ (.A(_00678_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _05496_ (.A0(net4091),
    .A1(_00185_),
    .S(_00677_),
    .X(_00679_));
 sky130_fd_sc_hd__clkbuf_1 _05497_ (.A(_00679_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _05498_ (.A0(net3997),
    .A1(_00189_),
    .S(_00677_),
    .X(_00680_));
 sky130_fd_sc_hd__clkbuf_1 _05499_ (.A(_00680_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _05500_ (.A0(net3354),
    .A1(_00528_),
    .S(_00677_),
    .X(_00681_));
 sky130_fd_sc_hd__clkbuf_1 _05501_ (.A(_00681_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[15] ));
 sky130_fd_sc_hd__a41oi_4 _05502_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[4] ),
    .A2(_00657_),
    .A3(_00658_),
    .A4(_00660_),
    .B1(_00181_),
    .Y(_00682_));
 sky130_fd_sc_hd__mux2_1 _05503_ (.A0(_00540_),
    .A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[16] ),
    .S(_00682_),
    .X(_00683_));
 sky130_fd_sc_hd__clkbuf_1 _05504_ (.A(_00683_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[16] ));
 sky130_fd_sc_hd__mux2_1 _05505_ (.A0(_00549_),
    .A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[17] ),
    .S(_00682_),
    .X(_00684_));
 sky130_fd_sc_hd__clkbuf_1 _05506_ (.A(_00684_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[17] ));
 sky130_fd_sc_hd__mux2_1 _05507_ (.A0(_00552_),
    .A1(net3915),
    .S(_00682_),
    .X(_00685_));
 sky130_fd_sc_hd__clkbuf_1 _05508_ (.A(_00685_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[18] ));
 sky130_fd_sc_hd__mux2_1 _05509_ (.A0(_00297_),
    .A1(net3191),
    .S(_00682_),
    .X(_00686_));
 sky130_fd_sc_hd__clkbuf_1 _05510_ (.A(_00686_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41oi_4 _05511_ (.A1(net3041),
    .A2(_00657_),
    .A3(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[2] ),
    .A4(_00660_),
    .B1(_00181_),
    .Y(_00687_));
 sky130_fd_sc_hd__mux2_1 _05512_ (.A0(_00540_),
    .A1(net4047),
    .S(_00687_),
    .X(_00688_));
 sky130_fd_sc_hd__clkbuf_1 _05513_ (.A(_00688_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _05514_ (.A0(_00549_),
    .A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[21] ),
    .S(_00687_),
    .X(_00689_));
 sky130_fd_sc_hd__clkbuf_1 _05515_ (.A(_00689_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _05516_ (.A0(_00552_),
    .A1(net3142),
    .S(_00687_),
    .X(_00690_));
 sky130_fd_sc_hd__clkbuf_1 _05517_ (.A(_00690_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _05518_ (.A0(_00297_),
    .A1(net247),
    .S(_00687_),
    .X(_00691_));
 sky130_fd_sc_hd__clkbuf_1 _05519_ (.A(_00691_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[23] ));
 sky130_fd_sc_hd__buf_6 _05520_ (.A(_00235_),
    .X(_00692_));
 sky130_fd_sc_hd__a41o_2 _05521_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[4] ),
    .A2(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ),
    .A3(_00658_),
    .A4(_00660_),
    .B1(_00522_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _05522_ (.A0(net4007),
    .A1(_00692_),
    .S(_00693_),
    .X(_00694_));
 sky130_fd_sc_hd__clkbuf_1 _05523_ (.A(_00694_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[24] ));
 sky130_fd_sc_hd__buf_6 _05524_ (.A(_00292_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _05525_ (.A0(net4040),
    .A1(_00695_),
    .S(_00693_),
    .X(_00696_));
 sky130_fd_sc_hd__clkbuf_1 _05526_ (.A(_00696_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[25] ));
 sky130_fd_sc_hd__buf_6 _05527_ (.A(_00188_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _05528_ (.A0(net4108),
    .A1(_00697_),
    .S(_00693_),
    .X(_00698_));
 sky130_fd_sc_hd__clkbuf_1 _05529_ (.A(_00698_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _05530_ (.A0(net3169),
    .A1(_00528_),
    .S(_00693_),
    .X(_00699_));
 sky130_fd_sc_hd__clkbuf_1 _05531_ (.A(_00699_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41oi_4 _05532_ (.A1(net3534),
    .A2(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ),
    .A3(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[2] ),
    .A4(_00660_),
    .B1(_00181_),
    .Y(_00700_));
 sky130_fd_sc_hd__mux2_1 _05533_ (.A0(_00540_),
    .A1(net3951),
    .S(_00700_),
    .X(_00701_));
 sky130_fd_sc_hd__clkbuf_1 _05534_ (.A(_00701_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _05535_ (.A0(_00549_),
    .A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[29] ),
    .S(_00700_),
    .X(_00702_));
 sky130_fd_sc_hd__clkbuf_1 _05536_ (.A(_00702_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _05537_ (.A0(_00552_),
    .A1(net4016),
    .S(_00700_),
    .X(_00703_));
 sky130_fd_sc_hd__clkbuf_1 _05538_ (.A(_00703_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _05539_ (.A0(_00297_),
    .A1(net3646),
    .S(_00700_),
    .X(_00704_));
 sky130_fd_sc_hd__clkbuf_1 _05540_ (.A(_00704_),
    .X(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _05541_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .Y(_00705_));
 sky130_fd_sc_hd__inv_2 _05542_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .Y(_00706_));
 sky130_fd_sc_hd__a31o_1 _05543_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .A2(_00706_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_00707_));
 sky130_fd_sc_hd__or3b_1 _05544_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .B(_00707_),
    .C_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .X(_00708_));
 sky130_fd_sc_hd__o21ai_1 _05545_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fds ),
    .A2(_00705_),
    .B1(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _05546_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .B(_00707_),
    .Y(_00710_));
 sky130_fd_sc_hd__mux4_1 _05547_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_00711_));
 sky130_fd_sc_hd__nor2_1 _05548_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .B(_00711_),
    .Y(_00712_));
 sky130_fd_sc_hd__mux2_1 _05549_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(_00713_));
 sky130_fd_sc_hd__nand2_1 _05550_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .B(_00713_),
    .Y(_00714_));
 sky130_fd_sc_hd__inv_2 _05551_ (.A(net3988),
    .Y(_00715_));
 sky130_fd_sc_hd__mux2_1 _05552_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(_00716_));
 sky130_fd_sc_hd__nand2_1 _05553_ (.A(_00715_),
    .B(_00716_),
    .Y(_00717_));
 sky130_fd_sc_hd__inv_2 _05554_ (.A(net3616),
    .Y(_00718_));
 sky130_fd_sc_hd__a31o_1 _05555_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .A2(_00714_),
    .A3(_00717_),
    .B1(_00718_),
    .X(_00719_));
 sky130_fd_sc_hd__mux4_1 _05556_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_00720_));
 sky130_fd_sc_hd__mux4_1 _05557_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_00721_));
 sky130_fd_sc_hd__inv_2 _05558_ (.A(net3809),
    .Y(_00722_));
 sky130_fd_sc_hd__mux2_1 _05559_ (.A0(_00720_),
    .A1(_00721_),
    .S(_00722_),
    .X(_00723_));
 sky130_fd_sc_hd__a2bb2o_1 _05560_ (.A1_N(_00712_),
    .A2_N(_00719_),
    .B1(_00723_),
    .B2(_00718_),
    .X(_00724_));
 sky130_fd_sc_hd__and2b_1 _05561_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .X(_00725_));
 sky130_fd_sc_hd__a21bo_1 _05562_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _05563_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .X(_00727_));
 sky130_fd_sc_hd__o221a_1 _05564_ (.A1(_00725_),
    .A2(_00726_),
    .B1(_00727_),
    .B2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .X(_00728_));
 sky130_fd_sc_hd__inv_2 _05565_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .Y(_00729_));
 sky130_fd_sc_hd__mux4_1 _05566_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_00730_));
 sky130_fd_sc_hd__a21bo_1 _05567_ (.A1(_00729_),
    .A2(_00730_),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(_00731_));
 sky130_fd_sc_hd__mux4_1 _05568_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_00732_));
 sky130_fd_sc_hd__mux4_1 _05569_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _05570_ (.A0(_00732_),
    .A1(_00733_),
    .S(_00729_),
    .X(_00734_));
 sky130_fd_sc_hd__o22a_4 _05571_ (.A1(_00728_),
    .A2(_00731_),
    .B1(_00734_),
    .B2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _05572_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ),
    .S(_00735_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _05573_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ),
    .S(_00735_),
    .X(_00737_));
 sky130_fd_sc_hd__mux4_1 _05574_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_00738_));
 sky130_fd_sc_hd__nor2_1 _05575_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .B(_00738_),
    .Y(_00739_));
 sky130_fd_sc_hd__mux2_1 _05576_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(_00740_));
 sky130_fd_sc_hd__nand2_1 _05577_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .B(_00740_),
    .Y(_00741_));
 sky130_fd_sc_hd__mux2_1 _05578_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(_00742_));
 sky130_fd_sc_hd__or2b_1 _05579_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .B_N(_00742_),
    .X(_00743_));
 sky130_fd_sc_hd__inv_2 _05580_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .Y(_00744_));
 sky130_fd_sc_hd__a31o_1 _05581_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .A2(_00741_),
    .A3(_00743_),
    .B1(_00744_),
    .X(_00745_));
 sky130_fd_sc_hd__mux4_1 _05582_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_00746_));
 sky130_fd_sc_hd__mux4_1 _05583_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _05584_ (.A0(_00746_),
    .A1(_00747_),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(_00748_));
 sky130_fd_sc_hd__a2bb2o_2 _05585_ (.A1_N(_00739_),
    .A2_N(_00745_),
    .B1(_00748_),
    .B2(_00744_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _05586_ (.A0(_00736_),
    .A1(_00737_),
    .S(_00749_),
    .X(_00750_));
 sky130_fd_sc_hd__and2b_1 _05587_ (.A_N(_00724_),
    .B(_00750_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _05588_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ),
    .S(_00735_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _05589_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ),
    .S(_00735_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _05590_ (.A0(_00752_),
    .A1(_00753_),
    .S(_00749_),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _05591_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _05592_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00756_));
 sky130_fd_sc_hd__or2b_1 _05593_ (.A(_00756_),
    .B_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .X(_00757_));
 sky130_fd_sc_hd__o211a_1 _05594_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_00755_),
    .B1(_00757_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _05595_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00759_));
 sky130_fd_sc_hd__and2b_1 _05596_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .X(_00760_));
 sky130_fd_sc_hd__a21bo_1 _05597_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .X(_00761_));
 sky130_fd_sc_hd__inv_2 _05598_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .Y(_00762_));
 sky130_fd_sc_hd__o221a_1 _05599_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_00759_),
    .B1(_00760_),
    .B2(_00761_),
    .C1(_00762_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _05600_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00764_));
 sky130_fd_sc_hd__or3b_1 _05601_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .C_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .X(_00765_));
 sky130_fd_sc_hd__o211a_1 _05602_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_00764_),
    .B1(_00765_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _05603_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00767_));
 sky130_fd_sc_hd__inv_2 _05604_ (.A(_00767_),
    .Y(_00768_));
 sky130_fd_sc_hd__mux2_1 _05605_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00769_));
 sky130_fd_sc_hd__nor2_1 _05606_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .B(_00769_),
    .Y(_00770_));
 sky130_fd_sc_hd__a211o_1 _05607_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_00768_),
    .B1(_00770_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_00771_));
 sky130_fd_sc_hd__nand2_1 _05608_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .B(_00771_),
    .Y(_00772_));
 sky130_fd_sc_hd__o32a_1 _05609_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .A2(_00758_),
    .A3(_00763_),
    .B1(_00766_),
    .B2(_00772_),
    .X(_00773_));
 sky130_fd_sc_hd__a21bo_1 _05610_ (.A1(_00724_),
    .A2(_00754_),
    .B1_N(_00773_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _05611_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ),
    .S(_00735_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _05612_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ),
    .S(_00735_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _05613_ (.A0(_00775_),
    .A1(_00776_),
    .S(_00749_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _05614_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ),
    .S(_00735_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _05615_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ),
    .S(_00735_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _05616_ (.A0(_00778_),
    .A1(_00779_),
    .S(_00749_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _05617_ (.A0(_00777_),
    .A1(_00780_),
    .S(_00724_),
    .X(_00781_));
 sky130_fd_sc_hd__inv_8 _05618_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ),
    .Y(_00782_));
 sky130_fd_sc_hd__o221ai_4 _05619_ (.A1(_00751_),
    .A2(_00774_),
    .B1(_00781_),
    .B2(_00773_),
    .C1(_00782_),
    .Y(_00783_));
 sky130_fd_sc_hd__a22o_4 _05620_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .A2(_00709_),
    .B1(_00710_),
    .B2(_00783_),
    .X(_00784_));
 sky130_fd_sc_hd__inv_2 _05621_ (.A(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hd__clkbuf_4 _05622_ (.A(_00785_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__inv_2 _05623_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .Y(_00786_));
 sky130_fd_sc_hd__inv_2 _05624_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ),
    .Y(_00787_));
 sky130_fd_sc_hd__buf_2 _05625_ (.A(_00787_),
    .X(_00788_));
 sky130_fd_sc_hd__inv_2 _05626_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .Y(_00789_));
 sky130_fd_sc_hd__mux4_1 _05627_ (.A0(_00784_),
    .A1(_00786_),
    .A2(_00788_),
    .A3(_00789_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .X(_00790_));
 sky130_fd_sc_hd__clkinv_2 _05628_ (.A(_00790_),
    .Y(_00791_));
 sky130_fd_sc_hd__buf_2 _05629_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .X(_00792_));
 sky130_fd_sc_hd__buf_2 _05630_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .X(_00793_));
 sky130_fd_sc_hd__mux4_1 _05631_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(_00792_),
    .A3(_00793_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _05632_ (.A0(_00791_),
    .A1(_00794_),
    .S(net3171),
    .X(_00795_));
 sky130_fd_sc_hd__clkbuf_1 _05633_ (.A(net3172),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ));
 sky130_fd_sc_hd__inv_2 _05634_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .Y(_00796_));
 sky130_fd_sc_hd__a31o_1 _05635_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .A2(_00796_),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_00797_));
 sky130_fd_sc_hd__nand2_1 _05636_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .B(_00797_),
    .Y(_00798_));
 sky130_fd_sc_hd__inv_2 _05637_ (.A(net3659),
    .Y(_00799_));
 sky130_fd_sc_hd__mux4_1 _05638_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_00800_));
 sky130_fd_sc_hd__mux4_1 _05639_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _05640_ (.A0(_00800_),
    .A1(_00801_),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .X(_00802_));
 sky130_fd_sc_hd__mux4_1 _05641_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_00803_));
 sky130_fd_sc_hd__inv_2 _05642_ (.A(net3869),
    .Y(_00804_));
 sky130_fd_sc_hd__inv_2 _05643_ (.A(net3953),
    .Y(_00805_));
 sky130_fd_sc_hd__or2_1 _05644_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(_00806_));
 sky130_fd_sc_hd__o211a_1 _05645_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .A2(_00804_),
    .B1(_00805_),
    .C1(_00806_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _05646_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(_00808_));
 sky130_fd_sc_hd__a21bo_1 _05647_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .A2(_00808_),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .X(_00809_));
 sky130_fd_sc_hd__o221a_1 _05648_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .A2(_00803_),
    .B1(_00807_),
    .B2(_00809_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ),
    .X(_00810_));
 sky130_fd_sc_hd__a21oi_2 _05649_ (.A1(_00799_),
    .A2(_00802_),
    .B1(_00810_),
    .Y(_00811_));
 sky130_fd_sc_hd__inv_2 _05650_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .Y(_00812_));
 sky130_fd_sc_hd__inv_2 _05651_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .Y(_00813_));
 sky130_fd_sc_hd__mux4_1 _05652_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_00814_));
 sky130_fd_sc_hd__and2_1 _05653_ (.A(_00813_),
    .B(_00814_),
    .X(_00815_));
 sky130_fd_sc_hd__and2b_1 _05654_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .X(_00816_));
 sky130_fd_sc_hd__a21bo_1 _05655_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _05656_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .X(_00818_));
 sky130_fd_sc_hd__o221a_1 _05657_ (.A1(_00816_),
    .A2(_00817_),
    .B1(_00818_),
    .B2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .X(_00819_));
 sky130_fd_sc_hd__mux4_1 _05658_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_00820_));
 sky130_fd_sc_hd__and2_1 _05659_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .B(_00820_),
    .X(_00821_));
 sky130_fd_sc_hd__mux4_1 _05660_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_00822_));
 sky130_fd_sc_hd__a21o_1 _05661_ (.A1(_00813_),
    .A2(_00822_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(_00823_));
 sky130_fd_sc_hd__o32a_4 _05662_ (.A1(_00812_),
    .A2(_00815_),
    .A3(_00819_),
    .B1(_00821_),
    .B2(_00823_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _05663_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ),
    .S(_00824_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _05664_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ),
    .S(_00824_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _05665_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(_00827_));
 sky130_fd_sc_hd__inv_2 _05666_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .Y(_00828_));
 sky130_fd_sc_hd__mux2_1 _05667_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(_00829_));
 sky130_fd_sc_hd__a21bo_1 _05668_ (.A1(_00828_),
    .A2(_00829_),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(_00830_));
 sky130_fd_sc_hd__a21o_1 _05669_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .A2(_00827_),
    .B1(_00830_),
    .X(_00831_));
 sky130_fd_sc_hd__mux4_1 _05670_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_00832_));
 sky130_fd_sc_hd__o21a_1 _05671_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .A2(_00832_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .X(_00833_));
 sky130_fd_sc_hd__mux4_1 _05672_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_00834_));
 sky130_fd_sc_hd__mux4_1 _05673_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _05674_ (.A0(_00834_),
    .A1(_00835_),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(_00836_));
 sky130_fd_sc_hd__inv_2 _05675_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .Y(_00837_));
 sky130_fd_sc_hd__a22o_2 _05676_ (.A1(_00831_),
    .A2(_00833_),
    .B1(_00836_),
    .B2(_00837_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _05677_ (.A0(_00825_),
    .A1(_00826_),
    .S(_00838_),
    .X(_00839_));
 sky130_fd_sc_hd__nand2_1 _05678_ (.A(_00811_),
    .B(_00839_),
    .Y(_00840_));
 sky130_fd_sc_hd__mux2_1 _05679_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _05680_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_00842_));
 sky130_fd_sc_hd__or2b_1 _05681_ (.A(_00842_),
    .B_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(_00843_));
 sky130_fd_sc_hd__o211a_1 _05682_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_00841_),
    .B1(_00843_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _05683_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_00845_));
 sky130_fd_sc_hd__and2b_1 _05684_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .X(_00846_));
 sky130_fd_sc_hd__a21bo_1 _05685_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(_00847_));
 sky130_fd_sc_hd__inv_2 _05686_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .Y(_00848_));
 sky130_fd_sc_hd__o221a_1 _05687_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_00845_),
    .B1(_00846_),
    .B2(_00847_),
    .C1(_00848_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _05688_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_00850_));
 sky130_fd_sc_hd__or3b_1 _05689_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .C_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(_00851_));
 sky130_fd_sc_hd__o211a_1 _05690_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_00850_),
    .B1(_00851_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _05691_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_00853_));
 sky130_fd_sc_hd__inv_2 _05692_ (.A(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__mux2_1 _05693_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_00855_));
 sky130_fd_sc_hd__nor2_1 _05694_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .B(_00855_),
    .Y(_00856_));
 sky130_fd_sc_hd__a211o_1 _05695_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_00854_),
    .B1(_00856_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_00857_));
 sky130_fd_sc_hd__nand2_1 _05696_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .B(_00857_),
    .Y(_00858_));
 sky130_fd_sc_hd__o32a_1 _05697_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .A2(_00844_),
    .A3(_00849_),
    .B1(_00852_),
    .B2(_00858_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _05698_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ),
    .S(_00824_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _05699_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ),
    .S(_00824_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _05700_ (.A0(_00860_),
    .A1(_00861_),
    .S(_00838_),
    .X(_00862_));
 sky130_fd_sc_hd__or2b_1 _05701_ (.A(_00811_),
    .B_N(_00862_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _05702_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ),
    .S(_00824_),
    .X(_00864_));
 sky130_fd_sc_hd__or2_1 _05703_ (.A(_00838_),
    .B(_00864_),
    .X(_00865_));
 sky130_fd_sc_hd__clkinv_2 _05704_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ),
    .Y(_00866_));
 sky130_fd_sc_hd__clkinv_2 _05705_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ),
    .Y(_00867_));
 sky130_fd_sc_hd__mux2_1 _05706_ (.A0(_00866_),
    .A1(_00867_),
    .S(_00824_),
    .X(_00868_));
 sky130_fd_sc_hd__a21oi_1 _05707_ (.A1(_00838_),
    .A2(_00868_),
    .B1(_00811_),
    .Y(_00869_));
 sky130_fd_sc_hd__mux2_1 _05708_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ),
    .S(_00824_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _05709_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ),
    .S(_00824_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _05710_ (.A0(_00870_),
    .A1(_00871_),
    .S(_00838_),
    .X(_00872_));
 sky130_fd_sc_hd__a221oi_1 _05711_ (.A1(_00865_),
    .A2(_00869_),
    .B1(_00872_),
    .B2(_00811_),
    .C1(_00859_),
    .Y(_00873_));
 sky130_fd_sc_hd__a311o_1 _05712_ (.A1(_00840_),
    .A2(_00859_),
    .A3(_00863_),
    .B1(_00873_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ),
    .X(_00874_));
 sky130_fd_sc_hd__inv_2 _05713_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .Y(_00875_));
 sky130_fd_sc_hd__or3b_1 _05714_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .B(_00797_),
    .C_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .X(_00876_));
 sky130_fd_sc_hd__o21ai_1 _05715_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ),
    .A2(_00875_),
    .B1(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__and2_1 _05716_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .B(_00877_),
    .X(_00878_));
 sky130_fd_sc_hd__a21o_2 _05717_ (.A1(_00798_),
    .A2(_00874_),
    .B1(_00878_),
    .X(_00879_));
 sky130_fd_sc_hd__inv_2 _05718_ (.A(_00879_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__buf_4 _05719_ (.A(_00879_),
    .X(_00880_));
 sky130_fd_sc_hd__inv_2 _05720_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .Y(_00881_));
 sky130_fd_sc_hd__inv_2 _05721_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .Y(_00882_));
 sky130_fd_sc_hd__inv_2 _05722_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .Y(_00883_));
 sky130_fd_sc_hd__mux4_1 _05723_ (.A0(_00880_),
    .A1(_00881_),
    .A2(_00882_),
    .A3(_00883_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .X(_00884_));
 sky130_fd_sc_hd__clkinv_2 _05724_ (.A(_00884_),
    .Y(_00885_));
 sky130_fd_sc_hd__buf_2 _05725_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .X(_00886_));
 sky130_fd_sc_hd__buf_2 _05726_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .X(_00887_));
 sky130_fd_sc_hd__buf_2 _05727_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .X(_00888_));
 sky130_fd_sc_hd__buf_2 _05728_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .X(_00889_));
 sky130_fd_sc_hd__mux4_1 _05729_ (.A0(_00886_),
    .A1(_00887_),
    .A2(_00888_),
    .A3(_00889_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _05730_ (.A0(_00885_),
    .A1(_00890_),
    .S(net3706),
    .X(_00891_));
 sky130_fd_sc_hd__clkbuf_1 _05731_ (.A(_00891_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ));
 sky130_fd_sc_hd__a31o_1 _05732_ (.A1(_00796_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_00892_));
 sky130_fd_sc_hd__nand2_2 _05733_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .B(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__mux2_1 _05734_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00894_));
 sky130_fd_sc_hd__or3b_1 _05735_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .C_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .X(_00895_));
 sky130_fd_sc_hd__o211a_1 _05736_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_00894_),
    .B1(_00895_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _05737_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00897_));
 sky130_fd_sc_hd__inv_2 _05738_ (.A(_00897_),
    .Y(_00898_));
 sky130_fd_sc_hd__mux2_1 _05739_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00899_));
 sky130_fd_sc_hd__nor2_1 _05740_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .B(_00899_),
    .Y(_00900_));
 sky130_fd_sc_hd__a211o_1 _05741_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_00898_),
    .B1(_00900_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_00901_));
 sky130_fd_sc_hd__nand2_1 _05742_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .B(_00901_),
    .Y(_00902_));
 sky130_fd_sc_hd__mux2_1 _05743_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00903_));
 sky130_fd_sc_hd__or2_1 _05744_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .B(_00903_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _05745_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00905_));
 sky130_fd_sc_hd__or2b_1 _05746_ (.A(_00905_),
    .B_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _05747_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_00907_));
 sky130_fd_sc_hd__and2b_1 _05748_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .X(_00908_));
 sky130_fd_sc_hd__a21bo_1 _05749_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .X(_00909_));
 sky130_fd_sc_hd__inv_2 _05750_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .Y(_00910_));
 sky130_fd_sc_hd__o221a_1 _05751_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_00907_),
    .B1(_00908_),
    .B2(_00909_),
    .C1(_00910_),
    .X(_00911_));
 sky130_fd_sc_hd__a311o_1 _05752_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .A2(_00904_),
    .A3(_00906_),
    .B1(_00911_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .X(_00912_));
 sky130_fd_sc_hd__o21ai_2 _05753_ (.A1(_00896_),
    .A2(_00902_),
    .B1(_00912_),
    .Y(_00913_));
 sky130_fd_sc_hd__inv_2 _05754_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .Y(_00914_));
 sky130_fd_sc_hd__mux4_1 _05755_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_00915_));
 sky130_fd_sc_hd__and2b_1 _05756_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .B(_00915_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _05757_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .X(_00917_));
 sky130_fd_sc_hd__and2b_1 _05758_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .X(_00918_));
 sky130_fd_sc_hd__a21bo_1 _05759_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_00919_));
 sky130_fd_sc_hd__o221a_1 _05760_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .A2(_00917_),
    .B1(_00918_),
    .B2(_00919_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .X(_00920_));
 sky130_fd_sc_hd__mux4_1 _05761_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_00921_));
 sky130_fd_sc_hd__and2b_1 _05762_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .B(_00921_),
    .X(_00922_));
 sky130_fd_sc_hd__mux4_1 _05763_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_00923_));
 sky130_fd_sc_hd__a21o_1 _05764_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .A2(_00923_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(_00924_));
 sky130_fd_sc_hd__o32a_4 _05765_ (.A1(_00914_),
    .A2(_00916_),
    .A3(_00920_),
    .B1(_00922_),
    .B2(_00924_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _05766_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ),
    .S(_00925_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _05767_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ),
    .S(_00925_),
    .X(_00927_));
 sky130_fd_sc_hd__mux4_1 _05768_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_00928_));
 sky130_fd_sc_hd__nor2_1 _05769_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .B(_00928_),
    .Y(_00929_));
 sky130_fd_sc_hd__mux4_1 _05770_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_00930_));
 sky130_fd_sc_hd__and2b_1 _05771_ (.A_N(_00930_),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(_00931_));
 sky130_fd_sc_hd__mux4_1 _05772_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _05773_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(_00933_));
 sky130_fd_sc_hd__and2b_1 _05774_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .B(_00933_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _05775_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(_00935_));
 sky130_fd_sc_hd__a21bo_1 _05776_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .A2(_00935_),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(_00936_));
 sky130_fd_sc_hd__o221ai_1 _05777_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .A2(_00932_),
    .B1(_00934_),
    .B2(_00936_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .Y(_00937_));
 sky130_fd_sc_hd__o31a_2 _05778_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .A2(_00929_),
    .A3(_00931_),
    .B1(_00937_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _05779_ (.A0(_00926_),
    .A1(_00927_),
    .S(_00938_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _05780_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ),
    .S(_00925_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _05781_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ),
    .S(_00925_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _05782_ (.A0(_00940_),
    .A1(_00941_),
    .S(_00938_),
    .X(_00942_));
 sky130_fd_sc_hd__inv_2 _05783_ (.A(net3841),
    .Y(_00943_));
 sky130_fd_sc_hd__mux4_1 _05784_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_00944_));
 sky130_fd_sc_hd__mux4_1 _05785_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _05786_ (.A0(_00944_),
    .A1(_00945_),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .X(_00946_));
 sky130_fd_sc_hd__mux4_1 _05787_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_00947_));
 sky130_fd_sc_hd__inv_2 _05788_ (.A(net3912),
    .Y(_00948_));
 sky130_fd_sc_hd__or2_1 _05789_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(_00949_));
 sky130_fd_sc_hd__o211a_1 _05790_ (.A1(_00948_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.half_q ),
    .B1(_00949_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_00950_));
 sky130_fd_sc_hd__inv_2 _05791_ (.A(net3973),
    .Y(_00951_));
 sky130_fd_sc_hd__mux2_1 _05792_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(_00952_));
 sky130_fd_sc_hd__inv_2 _05793_ (.A(net3734),
    .Y(_00953_));
 sky130_fd_sc_hd__a21o_1 _05794_ (.A1(_00951_),
    .A2(_00952_),
    .B1(_00953_),
    .X(_00954_));
 sky130_fd_sc_hd__o221a_1 _05795_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .A2(_00947_),
    .B1(_00950_),
    .B2(_00954_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ),
    .X(_00955_));
 sky130_fd_sc_hd__a21oi_2 _05796_ (.A1(_00943_),
    .A2(_00946_),
    .B1(_00955_),
    .Y(_00956_));
 sky130_fd_sc_hd__mux2_1 _05797_ (.A0(_00939_),
    .A1(_00942_),
    .S(_00956_),
    .X(_00957_));
 sky130_fd_sc_hd__inv_2 _05798_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ),
    .Y(_00958_));
 sky130_fd_sc_hd__nand2_1 _05799_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ),
    .B(_00925_),
    .Y(_00959_));
 sky130_fd_sc_hd__o211ai_1 _05800_ (.A1(_00958_),
    .A2(_00925_),
    .B1(_00938_),
    .C1(_00959_),
    .Y(_00960_));
 sky130_fd_sc_hd__mux2_1 _05801_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ),
    .S(_00925_),
    .X(_00961_));
 sky130_fd_sc_hd__o21ba_1 _05802_ (.A1(_00938_),
    .A2(_00961_),
    .B1_N(_00956_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _05803_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ),
    .S(_00925_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _05804_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ),
    .S(_00925_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _05805_ (.A0(_00963_),
    .A1(_00964_),
    .S(_00938_),
    .X(_00965_));
 sky130_fd_sc_hd__o21a_1 _05806_ (.A1(_00896_),
    .A2(_00902_),
    .B1(_00912_),
    .X(_00966_));
 sky130_fd_sc_hd__a221o_1 _05807_ (.A1(_00960_),
    .A2(_00962_),
    .B1(_00965_),
    .B2(_00956_),
    .C1(_00966_),
    .X(_00967_));
 sky130_fd_sc_hd__o211ai_4 _05808_ (.A1(_00913_),
    .A2(_00957_),
    .B1(_00967_),
    .C1(_00782_),
    .Y(_00968_));
 sky130_fd_sc_hd__or3b_1 _05809_ (.A(_00892_),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .X(_00969_));
 sky130_fd_sc_hd__o21ai_1 _05810_ (.A1(_00875_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ),
    .B1(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__and2_2 _05811_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .B(_00970_),
    .X(_00971_));
 sky130_fd_sc_hd__a21o_4 _05812_ (.A1(_00893_),
    .A2(_00968_),
    .B1(_00971_),
    .X(_00972_));
 sky130_fd_sc_hd__inv_6 _05813_ (.A(_00972_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__buf_2 _05814_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ),
    .X(_00973_));
 sky130_fd_sc_hd__mux4_1 _05815_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(_00973_),
    .A2(_00886_),
    .A3(_00887_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ),
    .X(_00974_));
 sky130_fd_sc_hd__buf_2 _05816_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .X(_00975_));
 sky130_fd_sc_hd__buf_2 _05817_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .X(_00976_));
 sky130_fd_sc_hd__mux4_1 _05818_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00888_),
    .A3(_00889_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _05819_ (.A0(_00974_),
    .A1(_00977_),
    .S(net3515),
    .X(_00978_));
 sky130_fd_sc_hd__clkbuf_1 _05820_ (.A(_00978_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ));
 sky130_fd_sc_hd__a31o_1 _05821_ (.A1(_00706_),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_00979_));
 sky130_fd_sc_hd__or3b_1 _05822_ (.A(_00979_),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .X(_00980_));
 sky130_fd_sc_hd__o21ai_1 _05823_ (.A1(_00705_),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fds ),
    .B1(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__nand2_1 _05824_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .B(_00979_),
    .Y(_00982_));
 sky130_fd_sc_hd__mux2_1 _05825_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(_00983_));
 sky130_fd_sc_hd__inv_2 _05826_ (.A(net3482),
    .Y(_00984_));
 sky130_fd_sc_hd__mux2_1 _05827_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(_00985_));
 sky130_fd_sc_hd__inv_2 _05828_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .Y(_00986_));
 sky130_fd_sc_hd__a21o_1 _05829_ (.A1(_00984_),
    .A2(_00985_),
    .B1(_00986_),
    .X(_00987_));
 sky130_fd_sc_hd__a21o_1 _05830_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .A2(_00983_),
    .B1(_00987_),
    .X(_00988_));
 sky130_fd_sc_hd__mux4_1 _05831_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_00989_));
 sky130_fd_sc_hd__or2_1 _05832_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .B(_00989_),
    .X(_00990_));
 sky130_fd_sc_hd__mux4_1 _05833_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_00991_));
 sky130_fd_sc_hd__or2_1 _05834_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .B(_00991_),
    .X(_00992_));
 sky130_fd_sc_hd__mux4_1 _05835_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_00993_));
 sky130_fd_sc_hd__inv_2 _05836_ (.A(net3987),
    .Y(_00994_));
 sky130_fd_sc_hd__o21a_1 _05837_ (.A1(_00986_),
    .A2(_00993_),
    .B1(_00994_),
    .X(_00995_));
 sky130_fd_sc_hd__a32oi_4 _05838_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ),
    .A2(_00988_),
    .A3(_00990_),
    .B1(_00992_),
    .B2(_00995_),
    .Y(_00996_));
 sky130_fd_sc_hd__mux2_1 _05839_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .X(_00997_));
 sky130_fd_sc_hd__and2b_1 _05840_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .X(_00998_));
 sky130_fd_sc_hd__a21bo_1 _05841_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_00999_));
 sky130_fd_sc_hd__o221a_1 _05842_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .A2(_00997_),
    .B1(_00998_),
    .B2(_00999_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .X(_01000_));
 sky130_fd_sc_hd__inv_2 _05843_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .Y(_01001_));
 sky130_fd_sc_hd__mux4_1 _05844_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01002_));
 sky130_fd_sc_hd__a21bo_1 _05845_ (.A1(_01001_),
    .A2(_01002_),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .X(_01003_));
 sky130_fd_sc_hd__mux4_1 _05846_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01004_));
 sky130_fd_sc_hd__mux4_1 _05847_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _05848_ (.A0(_01004_),
    .A1(_01005_),
    .S(_01001_),
    .X(_01006_));
 sky130_fd_sc_hd__o22a_4 _05849_ (.A1(_01000_),
    .A2(_01003_),
    .B1(_01006_),
    .B2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _05850_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ),
    .S(_01007_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _05851_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ),
    .S(_01007_),
    .X(_01009_));
 sky130_fd_sc_hd__inv_2 _05852_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .Y(_01010_));
 sky130_fd_sc_hd__mux4_1 _05853_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_01011_));
 sky130_fd_sc_hd__mux4_1 _05854_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _05855_ (.A0(_01011_),
    .A1(_01012_),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(_01013_));
 sky130_fd_sc_hd__mux4_1 _05856_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _05857_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(_01015_));
 sky130_fd_sc_hd__and2b_1 _05858_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .B(_01015_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _05859_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(_01017_));
 sky130_fd_sc_hd__a21bo_1 _05860_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .A2(_01017_),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(_01018_));
 sky130_fd_sc_hd__o221a_1 _05861_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .A2(_01014_),
    .B1(_01016_),
    .B2(_01018_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .X(_01019_));
 sky130_fd_sc_hd__a21oi_4 _05862_ (.A1(_01010_),
    .A2(_01013_),
    .B1(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__mux2_1 _05863_ (.A0(_01008_),
    .A1(_01009_),
    .S(_01020_),
    .X(_01021_));
 sky130_fd_sc_hd__nand2_1 _05864_ (.A(_00996_),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__a32o_1 _05865_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ),
    .A2(_00988_),
    .A3(_00990_),
    .B1(_00992_),
    .B2(_00995_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _05866_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ),
    .S(_01007_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _05867_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ),
    .S(_01007_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _05868_ (.A0(_01024_),
    .A1(_01025_),
    .S(_01020_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _05869_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01027_));
 sky130_fd_sc_hd__inv_2 _05870_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .Y(_01028_));
 sky130_fd_sc_hd__or3_1 _05871_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .C(_01028_),
    .X(_01029_));
 sky130_fd_sc_hd__o211ai_1 _05872_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01027_),
    .B1(_01029_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .Y(_01030_));
 sky130_fd_sc_hd__mux2_1 _05873_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _05874_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01032_));
 sky130_fd_sc_hd__o21ba_1 _05875_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01032_),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_01033_));
 sky130_fd_sc_hd__o21ai_1 _05876_ (.A1(_01028_),
    .A2(_01031_),
    .B1(_01033_),
    .Y(_01034_));
 sky130_fd_sc_hd__mux2_1 _05877_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01035_));
 sky130_fd_sc_hd__or2_1 _05878_ (.A(_01028_),
    .B(_01035_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _05879_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01037_));
 sky130_fd_sc_hd__o21a_1 _05880_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01037_),
    .B1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _05881_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _05882_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01040_));
 sky130_fd_sc_hd__o21ba_1 _05883_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01040_),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_01041_));
 sky130_fd_sc_hd__o21a_1 _05884_ (.A1(_01028_),
    .A2(_01039_),
    .B1(_01041_),
    .X(_01042_));
 sky130_fd_sc_hd__a211oi_1 _05885_ (.A1(_01036_),
    .A2(_01038_),
    .B1(_01042_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .Y(_01043_));
 sky130_fd_sc_hd__a31o_1 _05886_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .A2(_01030_),
    .A3(_01034_),
    .B1(_01043_),
    .X(_01044_));
 sky130_fd_sc_hd__a21oi_1 _05887_ (.A1(_01023_),
    .A2(_01026_),
    .B1(_01044_),
    .Y(_01045_));
 sky130_fd_sc_hd__mux2_1 _05888_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ),
    .S(_01007_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _05889_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ),
    .S(_01007_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _05890_ (.A0(_01046_),
    .A1(_01047_),
    .S(_01020_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _05891_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ),
    .S(_01007_),
    .X(_01049_));
 sky130_fd_sc_hd__o21ai_1 _05892_ (.A1(_01020_),
    .A2(_01049_),
    .B1(_01023_),
    .Y(_01050_));
 sky130_fd_sc_hd__inv_2 _05893_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ),
    .Y(_01051_));
 sky130_fd_sc_hd__nand2_1 _05894_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ),
    .B(_01007_),
    .Y(_01052_));
 sky130_fd_sc_hd__o211a_1 _05895_ (.A1(_01051_),
    .A2(_01007_),
    .B1(_01020_),
    .C1(_01052_),
    .X(_01053_));
 sky130_fd_sc_hd__o2bb2a_1 _05896_ (.A1_N(_00996_),
    .A2_N(_01048_),
    .B1(_01050_),
    .B2(_01053_),
    .X(_01054_));
 sky130_fd_sc_hd__a221o_2 _05897_ (.A1(_01022_),
    .A2(_01045_),
    .B1(_01054_),
    .B2(_01044_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ),
    .X(_01055_));
 sky130_fd_sc_hd__a22o_4 _05898_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .A2(_00981_),
    .B1(_00982_),
    .B2(_01055_),
    .X(_01056_));
 sky130_fd_sc_hd__inv_2 _05899_ (.A(_01056_),
    .Y(_01057_));
 sky130_fd_sc_hd__clkbuf_4 _05900_ (.A(_01057_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__inv_2 _05901_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .Y(_01058_));
 sky130_fd_sc_hd__buf_2 _05902_ (.A(_01058_),
    .X(_01059_));
 sky130_fd_sc_hd__inv_2 _05903_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .Y(_01060_));
 sky130_fd_sc_hd__buf_2 _05904_ (.A(_01060_),
    .X(_01061_));
 sky130_fd_sc_hd__mux4_1 _05905_ (.A0(_01056_),
    .A1(_01059_),
    .A2(_00788_),
    .A3(_01061_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .X(_01062_));
 sky130_fd_sc_hd__clkinv_2 _05906_ (.A(_01062_),
    .Y(_01063_));
 sky130_fd_sc_hd__mux4_1 _05907_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A3(_00793_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _05908_ (.A0(_01063_),
    .A1(_01064_),
    .S(net3516),
    .X(_01065_));
 sky130_fd_sc_hd__clkbuf_1 _05909_ (.A(_01065_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ));
 sky130_fd_sc_hd__a31o_1 _05910_ (.A1(_00706_),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_01066_));
 sky130_fd_sc_hd__or3b_1 _05911_ (.A(_01066_),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .X(_01067_));
 sky130_fd_sc_hd__o21ai_1 _05912_ (.A1(_00705_),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fds ),
    .B1(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hd__nand2_1 _05913_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .B(_01066_),
    .Y(_01069_));
 sky130_fd_sc_hd__inv_2 _05914_ (.A(net3847),
    .Y(_01070_));
 sky130_fd_sc_hd__mux4_1 _05915_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01071_));
 sky130_fd_sc_hd__mux4_1 _05916_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _05917_ (.A0(_01071_),
    .A1(_01072_),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .X(_01073_));
 sky130_fd_sc_hd__mux4_1 _05918_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01074_));
 sky130_fd_sc_hd__inv_2 _05919_ (.A(net3956),
    .Y(_01075_));
 sky130_fd_sc_hd__or2_1 _05920_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(_01076_));
 sky130_fd_sc_hd__o211a_1 _05921_ (.A1(_01075_),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.half_q ),
    .B1(_01076_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01077_));
 sky130_fd_sc_hd__inv_2 _05922_ (.A(net4060),
    .Y(_01078_));
 sky130_fd_sc_hd__mux2_1 _05923_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(_01079_));
 sky130_fd_sc_hd__inv_2 _05924_ (.A(net3819),
    .Y(_01080_));
 sky130_fd_sc_hd__a21o_1 _05925_ (.A1(_01078_),
    .A2(_01079_),
    .B1(_01080_),
    .X(_01081_));
 sky130_fd_sc_hd__o221a_1 _05926_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .A2(_01074_),
    .B1(_01077_),
    .B2(_01081_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ),
    .X(_01082_));
 sky130_fd_sc_hd__a21o_1 _05927_ (.A1(_01070_),
    .A2(_01073_),
    .B1(_01082_),
    .X(_01083_));
 sky130_fd_sc_hd__inv_2 _05928_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .Y(_01084_));
 sky130_fd_sc_hd__mux4_1 _05929_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01085_));
 sky130_fd_sc_hd__nand2_1 _05930_ (.A(_01084_),
    .B(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__mux2_1 _05931_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .X(_01087_));
 sky130_fd_sc_hd__and2b_1 _05932_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .X(_01088_));
 sky130_fd_sc_hd__a21bo_1 _05933_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01089_));
 sky130_fd_sc_hd__o221ai_2 _05934_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .A2(_01087_),
    .B1(_01088_),
    .B2(_01089_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .Y(_01090_));
 sky130_fd_sc_hd__mux4_1 _05935_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01091_));
 sky130_fd_sc_hd__nand2_1 _05936_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .B(_01091_),
    .Y(_01092_));
 sky130_fd_sc_hd__mux4_1 _05937_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01093_));
 sky130_fd_sc_hd__a21oi_1 _05938_ (.A1(_01084_),
    .A2(_01093_),
    .B1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .Y(_01094_));
 sky130_fd_sc_hd__a32o_4 _05939_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .A2(_01086_),
    .A3(_01090_),
    .B1(_01092_),
    .B2(_01094_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _05940_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ),
    .S(_01095_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _05941_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ),
    .S(_01095_),
    .X(_01097_));
 sky130_fd_sc_hd__mux4_1 _05942_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_01098_));
 sky130_fd_sc_hd__nor2_1 _05943_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .B(_01098_),
    .Y(_01099_));
 sky130_fd_sc_hd__mux2_1 _05944_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(_01100_));
 sky130_fd_sc_hd__nand2_1 _05945_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .B(_01100_),
    .Y(_01101_));
 sky130_fd_sc_hd__mux2_1 _05946_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(_01102_));
 sky130_fd_sc_hd__or2b_1 _05947_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .B_N(_01102_),
    .X(_01103_));
 sky130_fd_sc_hd__inv_2 _05948_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .Y(_01104_));
 sky130_fd_sc_hd__a31o_1 _05949_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .A2(_01101_),
    .A3(_01103_),
    .B1(_01104_),
    .X(_01105_));
 sky130_fd_sc_hd__mux4_1 _05950_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_01106_));
 sky130_fd_sc_hd__mux4_1 _05951_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _05952_ (.A0(_01106_),
    .A1(_01107_),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(_01108_));
 sky130_fd_sc_hd__a2bb2o_2 _05953_ (.A1_N(_01099_),
    .A2_N(_01105_),
    .B1(_01108_),
    .B2(_01104_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _05954_ (.A0(_01096_),
    .A1(_01097_),
    .S(_01109_),
    .X(_01110_));
 sky130_fd_sc_hd__and2b_1 _05955_ (.A_N(_01083_),
    .B(_01110_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _05956_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ),
    .S(_01095_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _05957_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ),
    .S(_01095_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _05958_ (.A0(_01112_),
    .A1(_01113_),
    .S(_01109_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _05959_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _05960_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01116_));
 sky130_fd_sc_hd__or2b_1 _05961_ (.A(_01116_),
    .B_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .X(_01117_));
 sky130_fd_sc_hd__o211a_1 _05962_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_01115_),
    .B1(_01117_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _05963_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01119_));
 sky130_fd_sc_hd__and2b_1 _05964_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .X(_01120_));
 sky130_fd_sc_hd__a21bo_1 _05965_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .X(_01121_));
 sky130_fd_sc_hd__inv_2 _05966_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .Y(_01122_));
 sky130_fd_sc_hd__o221a_1 _05967_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_01119_),
    .B1(_01120_),
    .B2(_01121_),
    .C1(_01122_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _05968_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01124_));
 sky130_fd_sc_hd__or3b_1 _05969_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .C_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .X(_01125_));
 sky130_fd_sc_hd__o211a_1 _05970_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_01124_),
    .B1(_01125_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _05971_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01127_));
 sky130_fd_sc_hd__inv_2 _05972_ (.A(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__mux2_1 _05973_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01129_));
 sky130_fd_sc_hd__nor2_1 _05974_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .B(_01129_),
    .Y(_01130_));
 sky130_fd_sc_hd__a211o_1 _05975_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_01128_),
    .B1(_01130_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(_01131_));
 sky130_fd_sc_hd__nand2_1 _05976_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .B(_01131_),
    .Y(_01132_));
 sky130_fd_sc_hd__o32a_1 _05977_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .A2(_01118_),
    .A3(_01123_),
    .B1(_01126_),
    .B2(_01132_),
    .X(_01133_));
 sky130_fd_sc_hd__a21bo_1 _05978_ (.A1(_01083_),
    .A2(_01114_),
    .B1_N(_01133_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _05979_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ),
    .S(_01095_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _05980_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ),
    .S(_01095_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _05981_ (.A0(_01135_),
    .A1(_01136_),
    .S(_01109_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _05982_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ),
    .S(_01095_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _05983_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ),
    .S(_01095_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _05984_ (.A0(_01138_),
    .A1(_01139_),
    .S(_01109_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _05985_ (.A0(_01137_),
    .A1(_01140_),
    .S(_01083_),
    .X(_01141_));
 sky130_fd_sc_hd__o221ai_4 _05986_ (.A1(_01111_),
    .A2(_01134_),
    .B1(_01141_),
    .B2(_01133_),
    .C1(_00782_),
    .Y(_01142_));
 sky130_fd_sc_hd__a22o_4 _05987_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .A2(_01068_),
    .B1(_01069_),
    .B2(_01142_),
    .X(_01143_));
 sky130_fd_sc_hd__inv_2 _05988_ (.A(_01143_),
    .Y(_01144_));
 sky130_fd_sc_hd__clkbuf_4 _05989_ (.A(_01144_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__mux4_1 _05990_ (.A0(_01143_),
    .A1(_01059_),
    .A2(_00788_),
    .A3(_01061_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .X(_01145_));
 sky130_fd_sc_hd__clkinv_2 _05991_ (.A(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__mux4_1 _05992_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A3(_00793_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _05993_ (.A0(_01146_),
    .A1(_01147_),
    .S(net3140),
    .X(_01148_));
 sky130_fd_sc_hd__clkbuf_1 _05994_ (.A(net3141),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ));
 sky130_fd_sc_hd__a31o_1 _05995_ (.A1(_00706_),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_01149_));
 sky130_fd_sc_hd__or3b_1 _05996_ (.A(_01149_),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .X(_01150_));
 sky130_fd_sc_hd__o21ai_1 _05997_ (.A1(_00705_),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fds ),
    .B1(_01150_),
    .Y(_01151_));
 sky130_fd_sc_hd__nand2_1 _05998_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .B(_01149_),
    .Y(_01152_));
 sky130_fd_sc_hd__inv_2 _05999_ (.A(net3716),
    .Y(_01153_));
 sky130_fd_sc_hd__mux4_1 _06000_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_01154_));
 sky130_fd_sc_hd__mux4_1 _06001_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _06002_ (.A0(_01154_),
    .A1(_01155_),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .X(_01156_));
 sky130_fd_sc_hd__mux4_1 _06003_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_01157_));
 sky130_fd_sc_hd__nor2_1 _06004_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .B(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__mux2_1 _06005_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(_01159_));
 sky130_fd_sc_hd__nand2_1 _06006_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .B(_01159_),
    .Y(_01160_));
 sky130_fd_sc_hd__inv_2 _06007_ (.A(net4065),
    .Y(_01161_));
 sky130_fd_sc_hd__mux2_1 _06008_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(_01162_));
 sky130_fd_sc_hd__nand2_1 _06009_ (.A(_01161_),
    .B(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__a31o_1 _06010_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .A2(_01160_),
    .A3(_01163_),
    .B1(_01153_),
    .X(_01164_));
 sky130_fd_sc_hd__o2bb2a_2 _06011_ (.A1_N(_01153_),
    .A2_N(_01156_),
    .B1(_01158_),
    .B2(_01164_),
    .X(_01165_));
 sky130_fd_sc_hd__and2b_1 _06012_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .X(_01166_));
 sky130_fd_sc_hd__a21bo_1 _06013_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _06014_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .X(_01168_));
 sky130_fd_sc_hd__o221a_1 _06015_ (.A1(_01166_),
    .A2(_01167_),
    .B1(_01168_),
    .B2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .X(_01169_));
 sky130_fd_sc_hd__inv_2 _06016_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .Y(_01170_));
 sky130_fd_sc_hd__mux4_1 _06017_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_01171_));
 sky130_fd_sc_hd__a21bo_1 _06018_ (.A1(_01170_),
    .A2(_01171_),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(_01172_));
 sky130_fd_sc_hd__mux4_1 _06019_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_01173_));
 sky130_fd_sc_hd__mux4_1 _06020_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _06021_ (.A0(_01173_),
    .A1(_01174_),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .X(_01175_));
 sky130_fd_sc_hd__o22a_4 _06022_ (.A1(_01169_),
    .A2(_01172_),
    .B1(_01175_),
    .B2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _06023_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ),
    .S(_01176_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _06024_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ),
    .S(_01176_),
    .X(_01178_));
 sky130_fd_sc_hd__mux4_1 _06025_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_01179_));
 sky130_fd_sc_hd__nor2_1 _06026_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .B(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__mux2_1 _06027_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(_01181_));
 sky130_fd_sc_hd__nand2_1 _06028_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .B(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__mux2_1 _06029_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(_01183_));
 sky130_fd_sc_hd__or2b_1 _06030_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .B_N(_01183_),
    .X(_01184_));
 sky130_fd_sc_hd__inv_2 _06031_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .Y(_01185_));
 sky130_fd_sc_hd__a31o_1 _06032_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .A2(_01182_),
    .A3(_01184_),
    .B1(_01185_),
    .X(_01186_));
 sky130_fd_sc_hd__mux4_1 _06033_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_01187_));
 sky130_fd_sc_hd__mux4_1 _06034_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _06035_ (.A0(_01187_),
    .A1(_01188_),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(_01189_));
 sky130_fd_sc_hd__a2bb2o_2 _06036_ (.A1_N(_01180_),
    .A2_N(_01186_),
    .B1(_01189_),
    .B2(_01185_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _06037_ (.A0(_01177_),
    .A1(_01178_),
    .S(_01190_),
    .X(_01191_));
 sky130_fd_sc_hd__nand2_1 _06038_ (.A(_01165_),
    .B(_01191_),
    .Y(_01192_));
 sky130_fd_sc_hd__inv_2 _06039_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .Y(_01193_));
 sky130_fd_sc_hd__mux2_1 _06040_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01194_));
 sky130_fd_sc_hd__inv_2 _06041_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .Y(_01195_));
 sky130_fd_sc_hd__or3_1 _06042_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .C(_01195_),
    .X(_01196_));
 sky130_fd_sc_hd__o211a_1 _06043_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_01194_),
    .B1(_01196_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _06044_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _06045_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01199_));
 sky130_fd_sc_hd__o21ba_1 _06046_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_01199_),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_01200_));
 sky130_fd_sc_hd__o21a_1 _06047_ (.A1(_01195_),
    .A2(_01198_),
    .B1(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _06048_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01202_));
 sky130_fd_sc_hd__or2_1 _06049_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .B(_01202_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _06050_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01204_));
 sky130_fd_sc_hd__or2_1 _06051_ (.A(_01195_),
    .B(_01204_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _06052_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _06053_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01207_));
 sky130_fd_sc_hd__o21ba_1 _06054_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_01207_),
    .B1_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_01208_));
 sky130_fd_sc_hd__o21a_1 _06055_ (.A1(_01195_),
    .A2(_01206_),
    .B1(_01208_),
    .X(_01209_));
 sky130_fd_sc_hd__a311o_1 _06056_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .A2(_01203_),
    .A3(_01205_),
    .B1(_01209_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .X(_01210_));
 sky130_fd_sc_hd__o31a_1 _06057_ (.A1(_01193_),
    .A2(_01197_),
    .A3(_01201_),
    .B1(_01210_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _06058_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ),
    .S(_01176_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _06059_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ),
    .S(_01176_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _06060_ (.A0(_01212_),
    .A1(_01213_),
    .S(_01190_),
    .X(_01214_));
 sky130_fd_sc_hd__or2b_1 _06061_ (.A(_01165_),
    .B_N(_01214_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _06062_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ),
    .S(_01176_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _06063_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ),
    .S(_01176_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _06064_ (.A0(_01216_),
    .A1(_01217_),
    .S(_01190_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _06065_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ),
    .S(_01176_),
    .X(_01219_));
 sky130_fd_sc_hd__or2_1 _06066_ (.A(_01190_),
    .B(_01219_),
    .X(_01220_));
 sky130_fd_sc_hd__clkinv_2 _06067_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ),
    .Y(_01221_));
 sky130_fd_sc_hd__clkinv_2 _06068_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ),
    .Y(_01222_));
 sky130_fd_sc_hd__mux2_1 _06069_ (.A0(_01221_),
    .A1(_01222_),
    .S(_01176_),
    .X(_01223_));
 sky130_fd_sc_hd__a21oi_1 _06070_ (.A1(_01190_),
    .A2(_01223_),
    .B1(_01165_),
    .Y(_01224_));
 sky130_fd_sc_hd__a221oi_1 _06071_ (.A1(_01165_),
    .A2(_01218_),
    .B1(_01220_),
    .B2(_01224_),
    .C1(_01211_),
    .Y(_01225_));
 sky130_fd_sc_hd__a311o_2 _06072_ (.A1(_01192_),
    .A2(_01211_),
    .A3(_01215_),
    .B1(_01225_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ),
    .X(_01226_));
 sky130_fd_sc_hd__a22o_4 _06073_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .A2(_01151_),
    .B1(_01152_),
    .B2(_01226_),
    .X(_01227_));
 sky130_fd_sc_hd__inv_2 _06074_ (.A(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__clkbuf_4 _06075_ (.A(_01228_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__inv_2 _06076_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .Y(_01229_));
 sky130_fd_sc_hd__mux4_1 _06077_ (.A0(_01227_),
    .A1(_01229_),
    .A2(_01059_),
    .A3(_01061_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .X(_01230_));
 sky130_fd_sc_hd__clkinv_2 _06078_ (.A(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__mux4_1 _06079_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A2(_00792_),
    .A3(_00793_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _06080_ (.A0(_01231_),
    .A1(_01232_),
    .S(net3148),
    .X(_01233_));
 sky130_fd_sc_hd__clkbuf_1 _06081_ (.A(net3149),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ));
 sky130_fd_sc_hd__a31o_1 _06082_ (.A1(_00796_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_01234_));
 sky130_fd_sc_hd__or3b_1 _06083_ (.A(_01234_),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .X(_01235_));
 sky130_fd_sc_hd__o21ai_1 _06084_ (.A1(_00875_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ),
    .B1(_01235_),
    .Y(_01236_));
 sky130_fd_sc_hd__nand2_1 _06085_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .B(_01234_),
    .Y(_01237_));
 sky130_fd_sc_hd__inv_2 _06086_ (.A(net3641),
    .Y(_01238_));
 sky130_fd_sc_hd__mux4_1 _06087_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_01239_));
 sky130_fd_sc_hd__mux4_1 _06088_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _06089_ (.A0(_01239_),
    .A1(_01240_),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .X(_01241_));
 sky130_fd_sc_hd__mux4_1 _06090_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_01242_));
 sky130_fd_sc_hd__nor2_1 _06091_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .B(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__mux2_1 _06092_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(_01244_));
 sky130_fd_sc_hd__nand2_1 _06093_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .B(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__inv_2 _06094_ (.A(net4036),
    .Y(_01246_));
 sky130_fd_sc_hd__mux2_1 _06095_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(_01247_));
 sky130_fd_sc_hd__nand2_1 _06096_ (.A(_01246_),
    .B(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__a31o_1 _06097_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .A2(_01245_),
    .A3(_01248_),
    .B1(_01238_),
    .X(_01249_));
 sky130_fd_sc_hd__o2bb2a_1 _06098_ (.A1_N(_01238_),
    .A2_N(_01241_),
    .B1(_01243_),
    .B2(_01249_),
    .X(_01250_));
 sky130_fd_sc_hd__inv_2 _06099_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .Y(_01251_));
 sky130_fd_sc_hd__inv_2 _06100_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .Y(_01252_));
 sky130_fd_sc_hd__mux4_1 _06101_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01253_));
 sky130_fd_sc_hd__and2_1 _06102_ (.A(_01252_),
    .B(_01253_),
    .X(_01254_));
 sky130_fd_sc_hd__and2b_1 _06103_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .X(_01255_));
 sky130_fd_sc_hd__a21bo_1 _06104_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _06105_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .X(_01257_));
 sky130_fd_sc_hd__o221a_1 _06106_ (.A1(_01255_),
    .A2(_01256_),
    .B1(_01257_),
    .B2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .X(_01258_));
 sky130_fd_sc_hd__mux4_1 _06107_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01259_));
 sky130_fd_sc_hd__and2_1 _06108_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .B(_01259_),
    .X(_01260_));
 sky130_fd_sc_hd__mux4_1 _06109_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01261_));
 sky130_fd_sc_hd__a21o_1 _06110_ (.A1(_01252_),
    .A2(_01261_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .X(_01262_));
 sky130_fd_sc_hd__o32a_4 _06111_ (.A1(_01251_),
    .A2(_01254_),
    .A3(_01258_),
    .B1(_01260_),
    .B2(_01262_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _06112_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ),
    .S(_01263_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _06113_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ),
    .S(_01263_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _06114_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(_01266_));
 sky130_fd_sc_hd__inv_2 _06115_ (.A(_01266_),
    .Y(_01267_));
 sky130_fd_sc_hd__mux2_1 _06116_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(_01268_));
 sky130_fd_sc_hd__nand2_1 _06117_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .B(_01268_),
    .Y(_01269_));
 sky130_fd_sc_hd__o211a_1 _06118_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .A2(_01267_),
    .B1(_01269_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(_01270_));
 sky130_fd_sc_hd__mux4_1 _06119_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_01271_));
 sky130_fd_sc_hd__o21ai_1 _06120_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .A2(_01271_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .Y(_01272_));
 sky130_fd_sc_hd__mux4_1 _06121_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_01273_));
 sky130_fd_sc_hd__mux4_1 _06122_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _06123_ (.A0(_01273_),
    .A1(_01274_),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(_01275_));
 sky130_fd_sc_hd__clkinv_2 _06124_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .Y(_01276_));
 sky130_fd_sc_hd__a2bb2o_2 _06125_ (.A1_N(_01270_),
    .A2_N(_01272_),
    .B1(_01275_),
    .B2(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _06126_ (.A0(_01264_),
    .A1(_01265_),
    .S(_01277_),
    .X(_01278_));
 sky130_fd_sc_hd__and2b_1 _06127_ (.A_N(_01250_),
    .B(_01278_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _06128_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ),
    .S(_01263_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _06129_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ),
    .S(_01263_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _06130_ (.A0(_01280_),
    .A1(_01281_),
    .S(_01277_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _06131_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _06132_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01284_));
 sky130_fd_sc_hd__or2b_1 _06133_ (.A(_01284_),
    .B_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .X(_01285_));
 sky130_fd_sc_hd__o211a_1 _06134_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01283_),
    .B1(_01285_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _06135_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01287_));
 sky130_fd_sc_hd__and2b_1 _06136_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .X(_01288_));
 sky130_fd_sc_hd__a21bo_1 _06137_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .X(_01289_));
 sky130_fd_sc_hd__inv_2 _06138_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .Y(_01290_));
 sky130_fd_sc_hd__o221a_1 _06139_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01287_),
    .B1(_01288_),
    .B2(_01289_),
    .C1(_01290_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _06140_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01292_));
 sky130_fd_sc_hd__or3b_1 _06141_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .C_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .X(_01293_));
 sky130_fd_sc_hd__o211a_1 _06142_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01292_),
    .B1(_01293_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _06143_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01295_));
 sky130_fd_sc_hd__inv_2 _06144_ (.A(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hd__mux2_1 _06145_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01297_));
 sky130_fd_sc_hd__nor2_1 _06146_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .B(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__a211o_1 _06147_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01296_),
    .B1(_01298_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_01299_));
 sky130_fd_sc_hd__nand2_1 _06148_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .B(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__o32a_1 _06149_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .A2(_01286_),
    .A3(_01291_),
    .B1(_01294_),
    .B2(_01300_),
    .X(_01301_));
 sky130_fd_sc_hd__a21bo_1 _06150_ (.A1(_01250_),
    .A2(_01282_),
    .B1_N(_01301_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _06151_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ),
    .S(_01263_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _06152_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ),
    .S(_01263_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _06153_ (.A0(_01303_),
    .A1(_01304_),
    .S(_01277_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _06154_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ),
    .S(_01263_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _06155_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ),
    .S(_01263_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _06156_ (.A0(_01306_),
    .A1(_01307_),
    .S(_01277_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _06157_ (.A0(_01305_),
    .A1(_01308_),
    .S(_01250_),
    .X(_01309_));
 sky130_fd_sc_hd__o221ai_4 _06158_ (.A1(_01279_),
    .A2(_01302_),
    .B1(_01309_),
    .B2(_01301_),
    .C1(_00782_),
    .Y(_01310_));
 sky130_fd_sc_hd__a22o_2 _06159_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .A2(_01236_),
    .B1(_01237_),
    .B2(_01310_),
    .X(_01311_));
 sky130_fd_sc_hd__clkinv_2 _06160_ (.A(_01311_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__mux4_1 _06161_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A1(_00973_),
    .A2(_00975_),
    .A3(_00976_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .X(_01312_));
 sky130_fd_sc_hd__mux4_1 _06162_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(_00887_),
    .A2(_00888_),
    .A3(_00889_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _06163_ (.A0(_01312_),
    .A1(_01313_),
    .S(net3285),
    .X(_01314_));
 sky130_fd_sc_hd__clkbuf_1 _06164_ (.A(net3286),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ));
 sky130_fd_sc_hd__a31o_1 _06165_ (.A1(_00796_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_01315_));
 sky130_fd_sc_hd__or3b_1 _06166_ (.A(_01315_),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .X(_01316_));
 sky130_fd_sc_hd__o21ai_1 _06167_ (.A1(_00875_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ),
    .B1(_01316_),
    .Y(_01317_));
 sky130_fd_sc_hd__nand2_1 _06168_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .B(_01315_),
    .Y(_01318_));
 sky130_fd_sc_hd__mux2_1 _06169_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(_01319_));
 sky130_fd_sc_hd__inv_2 _06170_ (.A(net3794),
    .Y(_01320_));
 sky130_fd_sc_hd__inv_2 _06171_ (.A(net3944),
    .Y(_01321_));
 sky130_fd_sc_hd__or2_1 _06172_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(_01322_));
 sky130_fd_sc_hd__o211a_1 _06173_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .A2(_01320_),
    .B1(_01321_),
    .C1(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__inv_2 _06174_ (.A(net3856),
    .Y(_01324_));
 sky130_fd_sc_hd__a211o_1 _06175_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .A2(_01319_),
    .B1(_01323_),
    .C1(_01324_),
    .X(_01325_));
 sky130_fd_sc_hd__mux4_1 _06176_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01326_));
 sky130_fd_sc_hd__o21a_1 _06177_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .A2(_01326_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ),
    .X(_01327_));
 sky130_fd_sc_hd__mux4_1 _06178_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01328_));
 sky130_fd_sc_hd__mux4_1 _06179_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _06180_ (.A0(_01328_),
    .A1(_01329_),
    .S(_01324_),
    .X(_01330_));
 sky130_fd_sc_hd__inv_2 _06181_ (.A(net3462),
    .Y(_01331_));
 sky130_fd_sc_hd__a22o_1 _06182_ (.A1(_01325_),
    .A2(_01327_),
    .B1(_01330_),
    .B2(_01331_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _06183_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .X(_01333_));
 sky130_fd_sc_hd__and2b_1 _06184_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .X(_01334_));
 sky130_fd_sc_hd__a21bo_1 _06185_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01335_));
 sky130_fd_sc_hd__o221a_1 _06186_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .A2(_01333_),
    .B1(_01334_),
    .B2(_01335_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .X(_01336_));
 sky130_fd_sc_hd__inv_2 _06187_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .Y(_01337_));
 sky130_fd_sc_hd__mux4_1 _06188_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01338_));
 sky130_fd_sc_hd__a21bo_1 _06189_ (.A1(_01337_),
    .A2(_01338_),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .X(_01339_));
 sky130_fd_sc_hd__mux4_1 _06190_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01340_));
 sky130_fd_sc_hd__mux4_1 _06191_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _06192_ (.A0(_01340_),
    .A1(_01341_),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .X(_01342_));
 sky130_fd_sc_hd__o22a_4 _06193_ (.A1(_01336_),
    .A2(_01339_),
    .B1(_01342_),
    .B2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _06194_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ),
    .S(_01343_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _06195_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ),
    .S(_01343_),
    .X(_01345_));
 sky130_fd_sc_hd__mux4_1 _06196_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _06197_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(_01347_));
 sky130_fd_sc_hd__and2b_1 _06198_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .B(_01347_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _06199_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(_01349_));
 sky130_fd_sc_hd__a21bo_1 _06200_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .A2(_01349_),
    .B1_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(_01350_));
 sky130_fd_sc_hd__o221a_1 _06201_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .A2(_01346_),
    .B1(_01348_),
    .B2(_01350_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .X(_01351_));
 sky130_fd_sc_hd__mux4_1 _06202_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_01352_));
 sky130_fd_sc_hd__mux4_1 _06203_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _06204_ (.A0(_01352_),
    .A1(_01353_),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(_01354_));
 sky130_fd_sc_hd__and2b_1 _06205_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .B(_01354_),
    .X(_01355_));
 sky130_fd_sc_hd__nor2_2 _06206_ (.A(_01351_),
    .B(_01355_),
    .Y(_01356_));
 sky130_fd_sc_hd__mux2_1 _06207_ (.A0(_01344_),
    .A1(_01345_),
    .S(_01356_),
    .X(_01357_));
 sky130_fd_sc_hd__or2b_1 _06208_ (.A(_01332_),
    .B_N(_01357_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _06209_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ),
    .S(_01343_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _06210_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ),
    .S(_01343_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _06211_ (.A0(_01359_),
    .A1(_01360_),
    .S(_01356_),
    .X(_01361_));
 sky130_fd_sc_hd__inv_2 _06212_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .Y(_01362_));
 sky130_fd_sc_hd__mux2_1 _06213_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _06214_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01364_));
 sky130_fd_sc_hd__or2_1 _06215_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .B(_01364_),
    .X(_01365_));
 sky130_fd_sc_hd__o211a_1 _06216_ (.A1(_01362_),
    .A2(_01363_),
    .B1(_01365_),
    .C1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _06217_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _06218_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01368_));
 sky130_fd_sc_hd__or2_1 _06219_ (.A(_01362_),
    .B(_01368_),
    .X(_01369_));
 sky130_fd_sc_hd__inv_2 _06220_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .Y(_01370_));
 sky130_fd_sc_hd__o211a_1 _06221_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_01367_),
    .B1(_01369_),
    .C1(_01370_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _06222_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01372_));
 sky130_fd_sc_hd__or2_1 _06223_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .B(_01372_),
    .X(_01373_));
 sky130_fd_sc_hd__o311a_1 _06224_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .A3(_01362_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .C1(_01373_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _06225_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _06226_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01376_));
 sky130_fd_sc_hd__or2_1 _06227_ (.A(_01362_),
    .B(_01376_),
    .X(_01377_));
 sky130_fd_sc_hd__o211a_1 _06228_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_01375_),
    .B1(_01377_),
    .C1(_01370_),
    .X(_01378_));
 sky130_fd_sc_hd__or3b_1 _06229_ (.A(_01374_),
    .B(_01378_),
    .C_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .X(_01379_));
 sky130_fd_sc_hd__o31ai_2 _06230_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .A2(_01366_),
    .A3(_01371_),
    .B1(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__a21oi_1 _06231_ (.A1(_01332_),
    .A2(_01361_),
    .B1(_01380_),
    .Y(_01381_));
 sky130_fd_sc_hd__clkinv_2 _06232_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ),
    .Y(_01382_));
 sky130_fd_sc_hd__inv_2 _06233_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ),
    .Y(_01383_));
 sky130_fd_sc_hd__mux2_1 _06234_ (.A0(_01382_),
    .A1(_01383_),
    .S(_01343_),
    .X(_01384_));
 sky130_fd_sc_hd__clkinv_2 _06235_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ),
    .Y(_01385_));
 sky130_fd_sc_hd__clkinv_2 _06236_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ),
    .Y(_01386_));
 sky130_fd_sc_hd__mux2_1 _06237_ (.A0(_01385_),
    .A1(_01386_),
    .S(_01343_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _06238_ (.A0(_01384_),
    .A1(_01387_),
    .S(_01356_),
    .X(_01388_));
 sky130_fd_sc_hd__and2b_1 _06239_ (.A_N(_01343_),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ),
    .X(_01389_));
 sky130_fd_sc_hd__a211o_1 _06240_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ),
    .A2(_01343_),
    .B1(_01355_),
    .C1(_01351_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _06241_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ),
    .S(_01343_),
    .X(_01391_));
 sky130_fd_sc_hd__o221ai_1 _06242_ (.A1(_01389_),
    .A2(_01390_),
    .B1(_01391_),
    .B2(_01356_),
    .C1(_01332_),
    .Y(_01392_));
 sky130_fd_sc_hd__o211a_1 _06243_ (.A1(_01332_),
    .A2(_01388_),
    .B1(_01392_),
    .C1(_01380_),
    .X(_01393_));
 sky130_fd_sc_hd__a211o_1 _06244_ (.A1(_01358_),
    .A2(_01381_),
    .B1(_01393_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ),
    .X(_01394_));
 sky130_fd_sc_hd__a22o_4 _06245_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .A2(_01317_),
    .B1(_01318_),
    .B2(_01394_),
    .X(_01395_));
 sky130_fd_sc_hd__clkinv_2 _06246_ (.A(_01395_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__mux4_1 _06247_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A1(_00973_),
    .A2(_00975_),
    .A3(_00976_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ),
    .X(_01396_));
 sky130_fd_sc_hd__mux4_1 _06248_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A2(_00888_),
    .A3(_00889_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _06249_ (.A0(_01396_),
    .A1(_01397_),
    .S(net3384),
    .X(_01398_));
 sky130_fd_sc_hd__clkbuf_1 _06250_ (.A(_01398_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ));
 sky130_fd_sc_hd__mux4_1 _06251_ (.A0(_00880_),
    .A1(_00881_),
    .A2(_00882_),
    .A3(_00883_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .X(_01399_));
 sky130_fd_sc_hd__clkinv_2 _06252_ (.A(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__mux4_1 _06253_ (.A0(_00886_),
    .A1(_00887_),
    .A2(_00888_),
    .A3(_00889_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _06254_ (.A0(_01400_),
    .A1(_01401_),
    .S(net3602),
    .X(_01402_));
 sky130_fd_sc_hd__clkbuf_1 _06255_ (.A(_01402_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ));
 sky130_fd_sc_hd__mux4_1 _06256_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(_00973_),
    .A2(_00886_),
    .A3(_00887_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ),
    .X(_01403_));
 sky130_fd_sc_hd__mux4_1 _06257_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00888_),
    .A3(_00889_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _06258_ (.A0(_01403_),
    .A1(_01404_),
    .S(net3484),
    .X(_01405_));
 sky130_fd_sc_hd__clkbuf_1 _06259_ (.A(_01405_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ));
 sky130_fd_sc_hd__inv_2 _06260_ (.A(net3532),
    .Y(_01406_));
 sky130_fd_sc_hd__mux4_1 _06261_ (.A0(_00975_),
    .A1(_00976_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A3(_00973_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .S1(_01406_),
    .X(_01407_));
 sky130_fd_sc_hd__mux4_1 _06262_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(_00887_),
    .A2(_00888_),
    .A3(_00889_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _06263_ (.A0(_01407_),
    .A1(_01408_),
    .S(net3518),
    .X(_01409_));
 sky130_fd_sc_hd__clkbuf_1 _06264_ (.A(_01409_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ));
 sky130_fd_sc_hd__mux4_1 _06265_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(_00886_),
    .A2(_00888_),
    .A3(_00889_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ),
    .X(_01410_));
 sky130_fd_sc_hd__inv_2 _06266_ (.A(net3711),
    .Y(_01411_));
 sky130_fd_sc_hd__mux4_1 _06267_ (.A0(_00975_),
    .A1(_00976_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A3(_00973_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .S1(_01411_),
    .X(_01412_));
 sky130_fd_sc_hd__inv_2 _06268_ (.A(net3418),
    .Y(_01413_));
 sky130_fd_sc_hd__mux2_1 _06269_ (.A0(_01410_),
    .A1(_01412_),
    .S(_01413_),
    .X(_01414_));
 sky130_fd_sc_hd__clkbuf_1 _06270_ (.A(net3419),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ));
 sky130_fd_sc_hd__buf_8 _06271_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ),
    .X(_01415_));
 sky130_fd_sc_hd__nand3b_2 _06272_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .B(_01415_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.cfgd ),
    .Y(_01416_));
 sky130_fd_sc_hd__or3_1 _06273_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_01417_));
 sky130_fd_sc_hd__or2_2 _06274_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_01417_),
    .X(_01418_));
 sky130_fd_sc_hd__o21a_1 _06275_ (.A1(_01416_),
    .A2(_01418_),
    .B1(_00408_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _06276_ (.A0(_00540_),
    .A1(net3613),
    .S(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__clkbuf_1 _06277_ (.A(_01420_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _06278_ (.A0(_00549_),
    .A1(net3529),
    .S(_01419_),
    .X(_01421_));
 sky130_fd_sc_hd__clkbuf_1 _06279_ (.A(_01421_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _06280_ (.A0(_00552_),
    .A1(net3511),
    .S(_01419_),
    .X(_01422_));
 sky130_fd_sc_hd__clkbuf_1 _06281_ (.A(_01422_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__buf_4 _06282_ (.A(_00191_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _06283_ (.A0(_01423_),
    .A1(net3430),
    .S(_01419_),
    .X(_01424_));
 sky130_fd_sc_hd__clkbuf_1 _06284_ (.A(_01424_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _06285_ (.A(net4189),
    .X(_01425_));
 sky130_fd_sc_hd__clkbuf_2 _06286_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ),
    .X(_01426_));
 sky130_fd_sc_hd__inv_2 _06287_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .Y(_01427_));
 sky130_fd_sc_hd__or4_1 _06288_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_01426_),
    .C(_01427_),
    .D(_01416_),
    .X(_01428_));
 sky130_fd_sc_hd__o21a_1 _06289_ (.A1(_01425_),
    .A2(_01428_),
    .B1(_00408_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _06290_ (.A0(_00540_),
    .A1(net3556),
    .S(_01429_),
    .X(_01430_));
 sky130_fd_sc_hd__clkbuf_1 _06291_ (.A(_01430_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _06292_ (.A0(_00549_),
    .A1(net3204),
    .S(_01429_),
    .X(_01431_));
 sky130_fd_sc_hd__clkbuf_1 _06293_ (.A(_01431_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _06294_ (.A0(_00552_),
    .A1(net3773),
    .S(_01429_),
    .X(_01432_));
 sky130_fd_sc_hd__clkbuf_1 _06295_ (.A(_01432_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _06296_ (.A0(_01423_),
    .A1(net3360),
    .S(_01429_),
    .X(_01433_));
 sky130_fd_sc_hd__clkbuf_1 _06297_ (.A(_01433_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__and3b_1 _06298_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .B(_01415_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.cfgd ),
    .X(_01434_));
 sky130_fd_sc_hd__nand2_1 _06299_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_01417_),
    .Y(_01435_));
 sky130_fd_sc_hd__and2_1 _06300_ (.A(_01418_),
    .B(_01435_),
    .X(_01436_));
 sky130_fd_sc_hd__inv_2 _06301_ (.A(_01425_),
    .Y(_01437_));
 sky130_fd_sc_hd__or3_1 _06302_ (.A(_01426_),
    .B(_01437_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_01438_));
 sky130_fd_sc_hd__nand2_2 _06303_ (.A(_00170_),
    .B(_01418_),
    .Y(_01439_));
 sky130_fd_sc_hd__nor2_1 _06304_ (.A(_01438_),
    .B(_01439_),
    .Y(_01440_));
 sky130_fd_sc_hd__inv_2 _06305_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .Y(_01441_));
 sky130_fd_sc_hd__and3b_1 _06306_ (.A_N(_01438_),
    .B(_01441_),
    .C(_01434_),
    .X(_01442_));
 sky130_fd_sc_hd__inv_2 _06307_ (.A(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__a32o_1 _06308_ (.A1(_01434_),
    .A2(_01436_),
    .A3(_01440_),
    .B1(_01443_),
    .B2(net3766),
    .X(_01444_));
 sky130_fd_sc_hd__a21o_1 _06309_ (.A1(_00279_),
    .A2(_01444_),
    .B1(_00210_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__clkinv_2 _06310_ (.A(net3469),
    .Y(_01445_));
 sky130_fd_sc_hd__buf_8 _06311_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ),
    .X(_01446_));
 sky130_fd_sc_hd__nand2_2 _06312_ (.A(_01446_),
    .B(_01418_),
    .Y(_01447_));
 sky130_fd_sc_hd__mux2_1 _06313_ (.A0(_01445_),
    .A1(_01447_),
    .S(_01442_),
    .X(_01448_));
 sky130_fd_sc_hd__o21ai_1 _06314_ (.A1(_00646_),
    .A2(_01448_),
    .B1(_00508_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__and2_1 _06315_ (.A(_00187_),
    .B(_01418_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _06316_ (.A0(net3572),
    .A1(_01449_),
    .S(_01442_),
    .X(_01450_));
 sky130_fd_sc_hd__a21o_1 _06317_ (.A1(_00279_),
    .A2(_01450_),
    .B1(_00222_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__clkinv_2 _06318_ (.A(net3564),
    .Y(_01451_));
 sky130_fd_sc_hd__buf_8 _06319_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ),
    .X(_01452_));
 sky130_fd_sc_hd__nand2_1 _06320_ (.A(_01452_),
    .B(_01418_),
    .Y(_01453_));
 sky130_fd_sc_hd__mux2_1 _06321_ (.A0(_01451_),
    .A1(_01453_),
    .S(_01442_),
    .X(_01454_));
 sky130_fd_sc_hd__o21ai_1 _06322_ (.A1(_00646_),
    .A2(_01454_),
    .B1(_00621_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_1 _06323_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_01416_),
    .Y(_01455_));
 sky130_fd_sc_hd__and3b_1 _06324_ (.A_N(_01426_),
    .B(_01425_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_01456_));
 sky130_fd_sc_hd__a21oi_2 _06325_ (.A1(_01455_),
    .A2(_01456_),
    .B1(_00267_),
    .Y(_01457_));
 sky130_fd_sc_hd__mux2_1 _06326_ (.A0(_00540_),
    .A1(net3507),
    .S(_01457_),
    .X(_01458_));
 sky130_fd_sc_hd__clkbuf_1 _06327_ (.A(_01458_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _06328_ (.A0(_00549_),
    .A1(net3366),
    .S(_01457_),
    .X(_01459_));
 sky130_fd_sc_hd__clkbuf_1 _06329_ (.A(_01459_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _06330_ (.A0(_00552_),
    .A1(net3551),
    .S(_01457_),
    .X(_01460_));
 sky130_fd_sc_hd__clkbuf_1 _06331_ (.A(_01460_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _06332_ (.A0(_01423_),
    .A1(net3567),
    .S(_01457_),
    .X(_01461_));
 sky130_fd_sc_hd__clkbuf_1 _06333_ (.A(_01461_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4_1 _06334_ (.A(_01426_),
    .B(_01437_),
    .C(_01427_),
    .D(_01455_),
    .X(_01462_));
 sky130_fd_sc_hd__clkbuf_2 _06335_ (.A(_01462_),
    .X(_01463_));
 sky130_fd_sc_hd__nand2_1 _06336_ (.A(_01439_),
    .B(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hd__or2_1 _06337_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .B(_01463_),
    .X(_01465_));
 sky130_fd_sc_hd__a31o_1 _06338_ (.A1(_00599_),
    .A2(_01464_),
    .A3(_01465_),
    .B1(_00603_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _06339_ (.A(_01447_),
    .B(_01463_),
    .Y(_01466_));
 sky130_fd_sc_hd__or2_1 _06340_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .B(_01463_),
    .X(_01467_));
 sky130_fd_sc_hd__a31o_1 _06341_ (.A1(_00599_),
    .A2(_01466_),
    .A3(_01467_),
    .B1(_00487_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__or2b_1 _06342_ (.A(_01449_),
    .B_N(_01463_),
    .X(_01468_));
 sky130_fd_sc_hd__or2_1 _06343_ (.A(net4024),
    .B(_01463_),
    .X(_01469_));
 sky130_fd_sc_hd__a31o_1 _06344_ (.A1(_00599_),
    .A2(_01468_),
    .A3(_01469_),
    .B1(_00394_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _06345_ (.A(net3863),
    .B(_01463_),
    .Y(_01470_));
 sky130_fd_sc_hd__buf_6 _06346_ (.A(_00236_),
    .X(_01471_));
 sky130_fd_sc_hd__a211o_1 _06347_ (.A1(_01453_),
    .A2(_01463_),
    .B1(_01470_),
    .C1(_01471_),
    .X(_01472_));
 sky130_fd_sc_hd__nand2_1 _06348_ (.A(_00263_),
    .B(_01472_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _06349_ (.A1(_01426_),
    .A2(_01437_),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .A4(_01455_),
    .B1(_00522_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _06350_ (.A0(net4076),
    .A1(_00692_),
    .S(_01473_),
    .X(_01474_));
 sky130_fd_sc_hd__clkbuf_1 _06351_ (.A(_01474_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _06352_ (.A0(net4179),
    .A1(_00695_),
    .S(_01473_),
    .X(_01475_));
 sky130_fd_sc_hd__clkbuf_1 _06353_ (.A(_01475_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _06354_ (.A0(net4044),
    .A1(_00697_),
    .S(_01473_),
    .X(_01476_));
 sky130_fd_sc_hd__clkbuf_1 _06355_ (.A(_01476_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _06356_ (.A0(net3853),
    .A1(_00528_),
    .S(_01473_),
    .X(_01477_));
 sky130_fd_sc_hd__clkbuf_1 _06357_ (.A(_01477_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_2 _06358_ (.A(_01426_),
    .B(_01425_),
    .C(_01427_),
    .D(_01455_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _06359_ (.A0(_00804_),
    .A1(_01439_),
    .S(_01478_),
    .X(_01479_));
 sky130_fd_sc_hd__o21ai_1 _06360_ (.A1(_00646_),
    .A2(_01479_),
    .B1(_00614_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _06361_ (.A0(_00805_),
    .A1(_01447_),
    .S(_01478_),
    .X(_01480_));
 sky130_fd_sc_hd__buf_4 _06362_ (.A(_00305_),
    .X(_01481_));
 sky130_fd_sc_hd__o21ai_1 _06363_ (.A1(_00646_),
    .A2(_01480_),
    .B1(_01481_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _06364_ (.A0(net4121),
    .A1(_01449_),
    .S(_01478_),
    .X(_01482_));
 sky130_fd_sc_hd__a21o_1 _06365_ (.A1(_00279_),
    .A2(_01482_),
    .B1(_00222_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _06366_ (.A0(_00799_),
    .A1(_01453_),
    .S(_01478_),
    .X(_01483_));
 sky130_fd_sc_hd__o21ai_1 _06367_ (.A1(_00646_),
    .A2(_01483_),
    .B1(_00621_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _06368_ (.A1(_01426_),
    .A2(_01425_),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .A4(_01455_),
    .B1(_00522_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _06369_ (.A0(net4175),
    .A1(_00692_),
    .S(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__clkbuf_1 _06370_ (.A(_01485_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _06371_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A1(_00695_),
    .S(_01484_),
    .X(_01486_));
 sky130_fd_sc_hd__clkbuf_1 _06372_ (.A(_01486_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _06373_ (.A0(net3901),
    .A1(_00697_),
    .S(_01484_),
    .X(_01487_));
 sky130_fd_sc_hd__clkbuf_1 _06374_ (.A(_01487_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _06375_ (.A0(net3975),
    .A1(_00528_),
    .S(_01484_),
    .X(_01488_));
 sky130_fd_sc_hd__clkbuf_1 _06376_ (.A(_01488_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__buf_6 _06377_ (.A(_00407_),
    .X(_01489_));
 sky130_fd_sc_hd__o31a_2 _06378_ (.A1(_01441_),
    .A2(_01416_),
    .A3(_01417_),
    .B1(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _06379_ (.A0(_00540_),
    .A1(net3830),
    .S(_01490_),
    .X(_01491_));
 sky130_fd_sc_hd__clkbuf_1 _06380_ (.A(_01491_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _06381_ (.A0(_00549_),
    .A1(net3202),
    .S(_01490_),
    .X(_01492_));
 sky130_fd_sc_hd__clkbuf_1 _06382_ (.A(_01492_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _06383_ (.A0(_00552_),
    .A1(net3872),
    .S(_01490_),
    .X(_01493_));
 sky130_fd_sc_hd__clkbuf_1 _06384_ (.A(_01493_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _06385_ (.A0(_01423_),
    .A1(net3875),
    .S(_01490_),
    .X(_01494_));
 sky130_fd_sc_hd__clkbuf_1 _06386_ (.A(_01494_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__clkbuf_4 _06387_ (.A(_00171_),
    .X(_01495_));
 sky130_fd_sc_hd__or2_1 _06388_ (.A(_01416_),
    .B(_01436_),
    .X(_01496_));
 sky130_fd_sc_hd__buf_8 _06389_ (.A(_00194_),
    .X(_01497_));
 sky130_fd_sc_hd__o41a_2 _06390_ (.A1(_01426_),
    .A2(_01425_),
    .A3(_01427_),
    .A4(_01496_),
    .B1(_01497_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _06391_ (.A0(_01495_),
    .A1(net3817),
    .S(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__clkbuf_1 _06392_ (.A(_01499_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__clkbuf_4 _06393_ (.A(_00184_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _06394_ (.A0(_01500_),
    .A1(net3625),
    .S(_01498_),
    .X(_01501_));
 sky130_fd_sc_hd__clkbuf_1 _06395_ (.A(_01501_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__inv_2 _06396_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .Y(_01502_));
 sky130_fd_sc_hd__inv_2 _06397_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .Y(_01503_));
 sky130_fd_sc_hd__a31o_1 _06398_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .A2(_01503_),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_01504_));
 sky130_fd_sc_hd__or3b_1 _06399_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .B(_01504_),
    .C_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .X(_01505_));
 sky130_fd_sc_hd__o21ai_1 _06400_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ),
    .A2(_01502_),
    .B1(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__nand2_1 _06401_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .B(_01504_),
    .Y(_01507_));
 sky130_fd_sc_hd__inv_2 _06402_ (.A(net3769),
    .Y(_01508_));
 sky130_fd_sc_hd__mux4_1 _06403_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_01509_));
 sky130_fd_sc_hd__mux4_1 _06404_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _06405_ (.A0(_01509_),
    .A1(_01510_),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .X(_01511_));
 sky130_fd_sc_hd__mux4_1 _06406_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_01512_));
 sky130_fd_sc_hd__inv_2 _06407_ (.A(net4022),
    .Y(_01513_));
 sky130_fd_sc_hd__or2_1 _06408_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(_01514_));
 sky130_fd_sc_hd__o211a_1 _06409_ (.A1(_01513_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.half_q ),
    .B1(_01514_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_01515_));
 sky130_fd_sc_hd__inv_2 _06410_ (.A(net3886),
    .Y(_01516_));
 sky130_fd_sc_hd__mux2_1 _06411_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(_01517_));
 sky130_fd_sc_hd__inv_2 _06412_ (.A(net3608),
    .Y(_01518_));
 sky130_fd_sc_hd__a21o_1 _06413_ (.A1(_01516_),
    .A2(_01517_),
    .B1(_01518_),
    .X(_01519_));
 sky130_fd_sc_hd__o221a_1 _06414_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .A2(_01512_),
    .B1(_01515_),
    .B2(_01519_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ),
    .X(_01520_));
 sky130_fd_sc_hd__a21o_1 _06415_ (.A1(_01508_),
    .A2(_01511_),
    .B1(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__and2b_1 _06416_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .X(_01522_));
 sky130_fd_sc_hd__a21bo_1 _06417_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _06418_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .X(_01524_));
 sky130_fd_sc_hd__o221a_1 _06419_ (.A1(_01522_),
    .A2(_01523_),
    .B1(_01524_),
    .B2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .X(_01525_));
 sky130_fd_sc_hd__inv_2 _06420_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .Y(_01526_));
 sky130_fd_sc_hd__mux4_1 _06421_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_01527_));
 sky130_fd_sc_hd__a21bo_1 _06422_ (.A1(_01526_),
    .A2(_01527_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(_01528_));
 sky130_fd_sc_hd__mux4_1 _06423_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_01529_));
 sky130_fd_sc_hd__mux4_1 _06424_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _06425_ (.A0(_01529_),
    .A1(_01530_),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .X(_01531_));
 sky130_fd_sc_hd__o22a_4 _06426_ (.A1(_01525_),
    .A2(_01528_),
    .B1(_01531_),
    .B2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _06427_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ),
    .S(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _06428_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ),
    .S(_01532_),
    .X(_01534_));
 sky130_fd_sc_hd__inv_2 _06429_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .Y(_01535_));
 sky130_fd_sc_hd__mux4_1 _06430_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_01536_));
 sky130_fd_sc_hd__mux4_1 _06431_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _06432_ (.A0(_01536_),
    .A1(_01537_),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(_01538_));
 sky130_fd_sc_hd__mux4_1 _06433_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _06434_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(_01540_));
 sky130_fd_sc_hd__and2b_1 _06435_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _06436_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(_01542_));
 sky130_fd_sc_hd__a21bo_1 _06437_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .A2(_01542_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(_01543_));
 sky130_fd_sc_hd__o221a_1 _06438_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .A2(_01539_),
    .B1(_01541_),
    .B2(_01543_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .X(_01544_));
 sky130_fd_sc_hd__a21oi_4 _06439_ (.A1(_01535_),
    .A2(_01538_),
    .B1(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__mux2_1 _06440_ (.A0(_01533_),
    .A1(_01534_),
    .S(_01545_),
    .X(_01546_));
 sky130_fd_sc_hd__and2b_1 _06441_ (.A_N(_01521_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _06442_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ),
    .S(_01532_),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _06443_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ),
    .S(_01532_),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _06444_ (.A0(_01548_),
    .A1(_01549_),
    .S(_01545_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _06445_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _06446_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01552_));
 sky130_fd_sc_hd__or2b_1 _06447_ (.A(_01552_),
    .B_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(_01553_));
 sky130_fd_sc_hd__o211a_1 _06448_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_01551_),
    .B1(_01553_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _06449_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01555_));
 sky130_fd_sc_hd__and2b_1 _06450_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .X(_01556_));
 sky130_fd_sc_hd__a21bo_1 _06451_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(_01557_));
 sky130_fd_sc_hd__inv_2 _06452_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .Y(_01558_));
 sky130_fd_sc_hd__o221a_1 _06453_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_01555_),
    .B1(_01556_),
    .B2(_01557_),
    .C1(_01558_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _06454_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01560_));
 sky130_fd_sc_hd__or3b_1 _06455_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .C_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(_01561_));
 sky130_fd_sc_hd__o211a_1 _06456_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_01560_),
    .B1(_01561_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _06457_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01563_));
 sky130_fd_sc_hd__inv_2 _06458_ (.A(_01563_),
    .Y(_01564_));
 sky130_fd_sc_hd__mux2_1 _06459_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_01565_));
 sky130_fd_sc_hd__nor2_1 _06460_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .B(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__a211o_1 _06461_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_01564_),
    .B1(_01566_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_01567_));
 sky130_fd_sc_hd__nand2_1 _06462_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__o32a_1 _06463_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .A2(_01554_),
    .A3(_01559_),
    .B1(_01562_),
    .B2(_01568_),
    .X(_01569_));
 sky130_fd_sc_hd__a21bo_1 _06464_ (.A1(_01521_),
    .A2(_01550_),
    .B1_N(_01569_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _06465_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ),
    .S(_01532_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _06466_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ),
    .S(_01532_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _06467_ (.A0(_01571_),
    .A1(_01572_),
    .S(_01545_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _06468_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ),
    .S(_01532_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _06469_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ),
    .S(_01532_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _06470_ (.A0(_01574_),
    .A1(_01575_),
    .S(_01545_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _06471_ (.A0(_01573_),
    .A1(_01576_),
    .S(_01521_),
    .X(_01577_));
 sky130_fd_sc_hd__buf_12 _06472_ (.A(_00782_),
    .X(_01578_));
 sky130_fd_sc_hd__o221ai_4 _06473_ (.A1(_01547_),
    .A2(_01570_),
    .B1(_01577_),
    .B2(_01569_),
    .C1(_01578_),
    .Y(_01579_));
 sky130_fd_sc_hd__a22o_4 _06474_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .A2(_01506_),
    .B1(_01507_),
    .B2(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__clkinv_2 _06475_ (.A(_01580_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__clkbuf_4 _06476_ (.A(_00551_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _06477_ (.A0(_01581_),
    .A1(net3799),
    .S(_01498_),
    .X(_01582_));
 sky130_fd_sc_hd__clkbuf_1 _06478_ (.A(_01582_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _06479_ (.A0(_01423_),
    .A1(net3386),
    .S(_01498_),
    .X(_01583_));
 sky130_fd_sc_hd__clkbuf_1 _06480_ (.A(_01583_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__buf_2 _06481_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .X(_01584_));
 sky130_fd_sc_hd__buf_2 _06482_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .X(_01585_));
 sky130_fd_sc_hd__mux4_1 _06483_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A2(_01584_),
    .A3(_01585_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .X(_01586_));
 sky130_fd_sc_hd__buf_2 _06484_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .X(_01587_));
 sky130_fd_sc_hd__buf_2 _06485_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .X(_01588_));
 sky130_fd_sc_hd__buf_2 _06486_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .X(_01589_));
 sky130_fd_sc_hd__buf_2 _06487_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .X(_01590_));
 sky130_fd_sc_hd__mux4_1 _06488_ (.A0(_01587_),
    .A1(_01588_),
    .A2(_01589_),
    .A3(_01590_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _06489_ (.A0(_01586_),
    .A1(_01591_),
    .S(net3157),
    .X(_01592_));
 sky130_fd_sc_hd__clkbuf_1 _06490_ (.A(_01592_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ));
 sky130_fd_sc_hd__nor2_2 _06491_ (.A(_01438_),
    .B(_01496_),
    .Y(_01593_));
 sky130_fd_sc_hd__or2_1 _06492_ (.A(net3791),
    .B(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__nand2_1 _06493_ (.A(_01439_),
    .B(_01593_),
    .Y(_01595_));
 sky130_fd_sc_hd__a31o_1 _06494_ (.A1(_00599_),
    .A2(_01594_),
    .A3(_01595_),
    .B1(_00603_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__a31o_1 _06495_ (.A1(_01503_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_01596_));
 sky130_fd_sc_hd__or3b_1 _06496_ (.A(_01596_),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .X(_01597_));
 sky130_fd_sc_hd__o21ai_1 _06497_ (.A1(_01502_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ),
    .B1(_01597_),
    .Y(_01598_));
 sky130_fd_sc_hd__nand2_1 _06498_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .B(_01596_),
    .Y(_01599_));
 sky130_fd_sc_hd__mux2_1 _06499_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_01600_));
 sky130_fd_sc_hd__inv_2 _06500_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .Y(_01601_));
 sky130_fd_sc_hd__or3_1 _06501_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .C(_01601_),
    .X(_01602_));
 sky130_fd_sc_hd__o211ai_1 _06502_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_01600_),
    .B1(_01602_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .Y(_01603_));
 sky130_fd_sc_hd__mux2_1 _06503_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_1 _06504_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_01605_));
 sky130_fd_sc_hd__o21ba_1 _06505_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_01605_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_01606_));
 sky130_fd_sc_hd__o21ai_1 _06506_ (.A1(_01601_),
    .A2(_01604_),
    .B1(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__mux2_1 _06507_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_01608_));
 sky130_fd_sc_hd__or2_1 _06508_ (.A(_01601_),
    .B(_01608_),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _06509_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_01610_));
 sky130_fd_sc_hd__o21a_1 _06510_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_01610_),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _06511_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _06512_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_01613_));
 sky130_fd_sc_hd__o21ba_1 _06513_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_01613_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_01614_));
 sky130_fd_sc_hd__o21a_1 _06514_ (.A1(_01601_),
    .A2(_01612_),
    .B1(_01614_),
    .X(_01615_));
 sky130_fd_sc_hd__a211oi_1 _06515_ (.A1(_01609_),
    .A2(_01611_),
    .B1(_01615_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .Y(_01616_));
 sky130_fd_sc_hd__a31o_1 _06516_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .A2(_01603_),
    .A3(_01607_),
    .B1(_01616_),
    .X(_01617_));
 sky130_fd_sc_hd__mux4_1 _06517_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_01618_));
 sky130_fd_sc_hd__or2_1 _06518_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .B(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _06519_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(_01620_));
 sky130_fd_sc_hd__inv_2 _06520_ (.A(net4035),
    .Y(_01621_));
 sky130_fd_sc_hd__mux2_1 _06521_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(_01622_));
 sky130_fd_sc_hd__inv_2 _06522_ (.A(net3905),
    .Y(_01623_));
 sky130_fd_sc_hd__a21o_1 _06523_ (.A1(_01621_),
    .A2(_01622_),
    .B1(_01623_),
    .X(_01624_));
 sky130_fd_sc_hd__a21o_1 _06524_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .A2(_01620_),
    .B1(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__mux4_1 _06525_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_01626_));
 sky130_fd_sc_hd__mux4_1 _06526_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_01627_));
 sky130_fd_sc_hd__or2_1 _06527_ (.A(_01623_),
    .B(_01627_),
    .X(_01628_));
 sky130_fd_sc_hd__inv_2 _06528_ (.A(net3938),
    .Y(_01629_));
 sky130_fd_sc_hd__o211a_1 _06529_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .A2(_01626_),
    .B1(_01628_),
    .C1(_01629_),
    .X(_01630_));
 sky130_fd_sc_hd__a31o_1 _06530_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ),
    .A2(_01619_),
    .A3(_01625_),
    .B1(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__and2b_1 _06531_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .X(_01632_));
 sky130_fd_sc_hd__a21bo_1 _06532_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _06533_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .X(_01634_));
 sky130_fd_sc_hd__o221a_1 _06534_ (.A1(_01632_),
    .A2(_01633_),
    .B1(_01634_),
    .B2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .X(_01635_));
 sky130_fd_sc_hd__inv_2 _06535_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .Y(_01636_));
 sky130_fd_sc_hd__mux4_1 _06536_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_01637_));
 sky130_fd_sc_hd__a21bo_1 _06537_ (.A1(_01636_),
    .A2(_01637_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(_01638_));
 sky130_fd_sc_hd__mux4_1 _06538_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_01639_));
 sky130_fd_sc_hd__mux4_1 _06539_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _06540_ (.A0(_01639_),
    .A1(_01640_),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .X(_01641_));
 sky130_fd_sc_hd__o22a_2 _06541_ (.A1(_01635_),
    .A2(_01638_),
    .B1(_01641_),
    .B2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _06542_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ),
    .S(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _06543_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ),
    .S(_01642_),
    .X(_01644_));
 sky130_fd_sc_hd__mux4_1 _06544_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _06545_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(_01646_));
 sky130_fd_sc_hd__and2b_1 _06546_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .B(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_1 _06547_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(_01648_));
 sky130_fd_sc_hd__a21bo_1 _06548_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .A2(_01648_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(_01649_));
 sky130_fd_sc_hd__o221a_1 _06549_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .A2(_01645_),
    .B1(_01647_),
    .B2(_01649_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .X(_01650_));
 sky130_fd_sc_hd__mux4_1 _06550_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_01651_));
 sky130_fd_sc_hd__mux4_1 _06551_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _06552_ (.A0(_01651_),
    .A1(_01652_),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(_01653_));
 sky130_fd_sc_hd__and2b_1 _06553_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .B(_01653_),
    .X(_01654_));
 sky130_fd_sc_hd__nor2_2 _06554_ (.A(_01650_),
    .B(_01654_),
    .Y(_01655_));
 sky130_fd_sc_hd__mux2_1 _06555_ (.A0(_01643_),
    .A1(_01644_),
    .S(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__nand2_1 _06556_ (.A(_01631_),
    .B(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__a31oi_2 _06557_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ),
    .A2(_01619_),
    .A3(_01625_),
    .B1(_01630_),
    .Y(_01658_));
 sky130_fd_sc_hd__mux2_1 _06558_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ),
    .S(_01642_),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _06559_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ),
    .S(_01642_),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _06560_ (.A0(_01659_),
    .A1(_01660_),
    .S(_01655_),
    .X(_01661_));
 sky130_fd_sc_hd__nand2_1 _06561_ (.A(_01658_),
    .B(_01661_),
    .Y(_01662_));
 sky130_fd_sc_hd__mux2_1 _06562_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ),
    .S(_01642_),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _06563_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ),
    .S(_01642_),
    .X(_01664_));
 sky130_fd_sc_hd__mux2_1 _06564_ (.A0(_01663_),
    .A1(_01664_),
    .S(_01655_),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _06565_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ),
    .S(_01642_),
    .X(_01666_));
 sky130_fd_sc_hd__o22ai_1 _06566_ (.A1(_01635_),
    .A2(_01638_),
    .B1(_01641_),
    .B2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .Y(_01667_));
 sky130_fd_sc_hd__o221a_1 _06567_ (.A1(_01635_),
    .A2(_01638_),
    .B1(_01641_),
    .B2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ),
    .X(_01668_));
 sky130_fd_sc_hd__a2111o_1 _06568_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ),
    .A2(_01667_),
    .B1(_01650_),
    .C1(_01654_),
    .D1(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__o211a_1 _06569_ (.A1(_01655_),
    .A2(_01666_),
    .B1(_01669_),
    .C1(_01658_),
    .X(_01670_));
 sky130_fd_sc_hd__a211oi_1 _06570_ (.A1(_01631_),
    .A2(_01665_),
    .B1(_01617_),
    .C1(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__a311o_2 _06571_ (.A1(_01617_),
    .A2(_01657_),
    .A3(_01662_),
    .B1(_01671_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ),
    .X(_01672_));
 sky130_fd_sc_hd__a22o_4 _06572_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .A2(_01598_),
    .B1(_01599_),
    .B2(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__clkinv_2 _06573_ (.A(_01673_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__nand2_1 _06574_ (.A(_01447_),
    .B(_01593_),
    .Y(_01674_));
 sky130_fd_sc_hd__or2_1 _06575_ (.A(net4130),
    .B(_01593_),
    .X(_01675_));
 sky130_fd_sc_hd__a31o_1 _06576_ (.A1(_00599_),
    .A2(_01674_),
    .A3(_01675_),
    .B1(_00487_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__buf_2 _06577_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ),
    .X(_01676_));
 sky130_fd_sc_hd__mux4_1 _06578_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(_01676_),
    .A2(_01587_),
    .A3(_01588_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(_01677_));
 sky130_fd_sc_hd__buf_2 _06579_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .X(_01678_));
 sky130_fd_sc_hd__mux4_1 _06580_ (.A0(_01678_),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(_01589_),
    .A3(_01590_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_1 _06581_ (.A0(_01677_),
    .A1(_01679_),
    .S(net3555),
    .X(_01680_));
 sky130_fd_sc_hd__clkbuf_1 _06582_ (.A(_01680_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ));
 sky130_fd_sc_hd__mux2_1 _06583_ (.A0(net3520),
    .A1(_01449_),
    .S(_01593_),
    .X(_01681_));
 sky130_fd_sc_hd__a21o_1 _06584_ (.A1(_00279_),
    .A2(_01681_),
    .B1(_00222_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__a31o_1 _06585_ (.A1(_01503_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_01682_));
 sky130_fd_sc_hd__or3b_1 _06586_ (.A(_01682_),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .X(_01683_));
 sky130_fd_sc_hd__o21ai_1 _06587_ (.A1(_01502_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ),
    .B1(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__nand2_1 _06588_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .B(_01682_),
    .Y(_01685_));
 sky130_fd_sc_hd__inv_2 _06589_ (.A(net3810),
    .Y(_01686_));
 sky130_fd_sc_hd__mux4_1 _06590_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_01687_));
 sky130_fd_sc_hd__mux4_1 _06591_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _06592_ (.A0(_01687_),
    .A1(_01688_),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .X(_01689_));
 sky130_fd_sc_hd__mux4_1 _06593_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_01690_));
 sky130_fd_sc_hd__inv_2 _06594_ (.A(net3885),
    .Y(_01691_));
 sky130_fd_sc_hd__inv_2 _06595_ (.A(net4127),
    .Y(_01692_));
 sky130_fd_sc_hd__or2_1 _06596_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(_01693_));
 sky130_fd_sc_hd__o211a_1 _06597_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .A2(_01691_),
    .B1(_01692_),
    .C1(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _06598_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(_01695_));
 sky130_fd_sc_hd__inv_2 _06599_ (.A(net3917),
    .Y(_01696_));
 sky130_fd_sc_hd__a21o_1 _06600_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .A2(_01695_),
    .B1(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__o221a_1 _06601_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .A2(_01690_),
    .B1(_01694_),
    .B2(_01697_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ),
    .X(_01698_));
 sky130_fd_sc_hd__a21oi_2 _06602_ (.A1(_01686_),
    .A2(_01689_),
    .B1(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__inv_2 _06603_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .Y(_01700_));
 sky130_fd_sc_hd__mux4_1 _06604_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01701_));
 sky130_fd_sc_hd__and2b_1 _06605_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .B(_01701_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _06606_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .X(_01703_));
 sky130_fd_sc_hd__and2b_1 _06607_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .X(_01704_));
 sky130_fd_sc_hd__a21bo_1 _06608_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01705_));
 sky130_fd_sc_hd__o221a_1 _06609_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .A2(_01703_),
    .B1(_01704_),
    .B2(_01705_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .X(_01706_));
 sky130_fd_sc_hd__mux4_1 _06610_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01707_));
 sky130_fd_sc_hd__and2b_1 _06611_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .B(_01707_),
    .X(_01708_));
 sky130_fd_sc_hd__mux4_1 _06612_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_01709_));
 sky130_fd_sc_hd__a21o_1 _06613_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .A2(_01709_),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .X(_01710_));
 sky130_fd_sc_hd__o32a_4 _06614_ (.A1(_01700_),
    .A2(_01702_),
    .A3(_01706_),
    .B1(_01708_),
    .B2(_01710_),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_1 _06615_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ),
    .S(_01711_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _06616_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ),
    .S(_01711_),
    .X(_01713_));
 sky130_fd_sc_hd__inv_2 _06617_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .Y(_01714_));
 sky130_fd_sc_hd__mux4_1 _06618_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_01715_));
 sky130_fd_sc_hd__mux4_1 _06619_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _06620_ (.A0(_01715_),
    .A1(_01716_),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(_01717_));
 sky130_fd_sc_hd__mux4_1 _06621_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_1 _06622_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(_01719_));
 sky130_fd_sc_hd__and2b_1 _06623_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .B(_01719_),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _06624_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(_01721_));
 sky130_fd_sc_hd__a21bo_1 _06625_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .A2(_01721_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(_01722_));
 sky130_fd_sc_hd__o221a_1 _06626_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .A2(_01718_),
    .B1(_01720_),
    .B2(_01722_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .X(_01723_));
 sky130_fd_sc_hd__a21o_2 _06627_ (.A1(_01714_),
    .A2(_01717_),
    .B1(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _06628_ (.A0(_01712_),
    .A1(_01713_),
    .S(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__and2_1 _06629_ (.A(_01699_),
    .B(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__inv_2 _06630_ (.A(_01699_),
    .Y(_01727_));
 sky130_fd_sc_hd__mux2_1 _06631_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ),
    .S(_01711_),
    .X(_01728_));
 sky130_fd_sc_hd__mux2_1 _06632_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ),
    .S(_01711_),
    .X(_01729_));
 sky130_fd_sc_hd__mux2_1 _06633_ (.A0(_01728_),
    .A1(_01729_),
    .S(_01724_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _06634_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01731_));
 sky130_fd_sc_hd__mux2_1 _06635_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01732_));
 sky130_fd_sc_hd__or2b_1 _06636_ (.A(_01732_),
    .B_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .X(_01733_));
 sky130_fd_sc_hd__o211a_1 _06637_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01731_),
    .B1(_01733_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_01734_));
 sky130_fd_sc_hd__mux2_1 _06638_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01735_));
 sky130_fd_sc_hd__and2b_1 _06639_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .X(_01736_));
 sky130_fd_sc_hd__a21bo_1 _06640_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .X(_01737_));
 sky130_fd_sc_hd__inv_2 _06641_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .Y(_01738_));
 sky130_fd_sc_hd__o221a_1 _06642_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01735_),
    .B1(_01736_),
    .B2(_01737_),
    .C1(_01738_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _06643_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01740_));
 sky130_fd_sc_hd__or3b_1 _06644_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .C_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .X(_01741_));
 sky130_fd_sc_hd__o211a_1 _06645_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01740_),
    .B1(_01741_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_01742_));
 sky130_fd_sc_hd__mux2_1 _06646_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01743_));
 sky130_fd_sc_hd__inv_2 _06647_ (.A(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__mux2_1 _06648_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_01745_));
 sky130_fd_sc_hd__nor2_1 _06649_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .B(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__a211o_1 _06650_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_01744_),
    .B1(_01746_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_01747_));
 sky130_fd_sc_hd__nand2_1 _06651_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__o32a_1 _06652_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .A2(_01734_),
    .A3(_01739_),
    .B1(_01742_),
    .B2(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__a21bo_1 _06653_ (.A1(_01727_),
    .A2(_01730_),
    .B1_N(_01749_),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _06654_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ),
    .S(_01711_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _06655_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ),
    .S(_01711_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _06656_ (.A0(_01751_),
    .A1(_01752_),
    .S(_01724_),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _06657_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ),
    .S(_01711_),
    .X(_01754_));
 sky130_fd_sc_hd__mux2_1 _06658_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ),
    .S(_01711_),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _06659_ (.A0(_01754_),
    .A1(_01755_),
    .S(_01724_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _06660_ (.A0(_01753_),
    .A1(_01756_),
    .S(_01699_),
    .X(_01757_));
 sky130_fd_sc_hd__o221ai_4 _06661_ (.A1(_01726_),
    .A2(_01750_),
    .B1(_01757_),
    .B2(_01749_),
    .C1(_01578_),
    .Y(_01758_));
 sky130_fd_sc_hd__a22o_4 _06662_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .A2(_01684_),
    .B1(_01685_),
    .B2(_01758_),
    .X(_01759_));
 sky130_fd_sc_hd__clkinv_2 _06663_ (.A(_01759_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__nor2_1 _06664_ (.A(net3804),
    .B(_01593_),
    .Y(_01760_));
 sky130_fd_sc_hd__a211o_1 _06665_ (.A1(_01453_),
    .A2(_01593_),
    .B1(_01760_),
    .C1(_01471_),
    .X(_01761_));
 sky130_fd_sc_hd__nand2_1 _06666_ (.A(_00263_),
    .B(_01761_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__clkbuf_4 _06667_ (.A(_00235_),
    .X(_01762_));
 sky130_fd_sc_hd__and3_2 _06668_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_01434_),
    .C(_01456_),
    .X(_01763_));
 sky130_fd_sc_hd__buf_8 _06669_ (.A(_00181_),
    .X(_01764_));
 sky130_fd_sc_hd__nor2_1 _06670_ (.A(_01764_),
    .B(_01763_),
    .Y(_01765_));
 sky130_fd_sc_hd__buf_4 _06671_ (.A(_00208_),
    .X(_01766_));
 sky130_fd_sc_hd__a221o_1 _06672_ (.A1(_01762_),
    .A2(_01763_),
    .B1(_01765_),
    .B2(net3227),
    .C1(_01766_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__inv_2 _06673_ (.A(net3658),
    .Y(_01767_));
 sky130_fd_sc_hd__mux4_1 _06674_ (.A0(_01678_),
    .A1(_01585_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A3(_01676_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .S1(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__mux4_1 _06675_ (.A0(_01584_),
    .A1(_01588_),
    .A2(_01589_),
    .A3(_01590_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _06676_ (.A0(_01768_),
    .A1(_01769_),
    .S(net3459),
    .X(_01770_));
 sky130_fd_sc_hd__clkbuf_1 _06677_ (.A(_01770_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ));
 sky130_fd_sc_hd__clkbuf_4 _06678_ (.A(_00292_),
    .X(_01771_));
 sky130_fd_sc_hd__clkbuf_8 _06679_ (.A(_00215_),
    .X(_01772_));
 sky130_fd_sc_hd__a221o_1 _06680_ (.A1(_01771_),
    .A2(_01763_),
    .B1(_01765_),
    .B2(net3207),
    .C1(_01772_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a31o_1 _06681_ (.A1(_01503_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_01773_));
 sky130_fd_sc_hd__or3b_1 _06682_ (.A(_01773_),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .X(_01774_));
 sky130_fd_sc_hd__o21ai_1 _06683_ (.A1(_01502_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ),
    .B1(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__nand2_1 _06684_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .B(_01773_),
    .Y(_01776_));
 sky130_fd_sc_hd__mux2_1 _06685_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01777_));
 sky130_fd_sc_hd__inv_2 _06686_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .Y(_01778_));
 sky130_fd_sc_hd__or3_1 _06687_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .C(_01778_),
    .X(_01779_));
 sky130_fd_sc_hd__o211ai_1 _06688_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_01777_),
    .B1(_01779_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .Y(_01780_));
 sky130_fd_sc_hd__mux2_1 _06689_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _06690_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01782_));
 sky130_fd_sc_hd__o21ba_1 _06691_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_01782_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(_01783_));
 sky130_fd_sc_hd__o21ai_1 _06692_ (.A1(_01778_),
    .A2(_01781_),
    .B1(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__mux2_1 _06693_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01785_));
 sky130_fd_sc_hd__or2_1 _06694_ (.A(_01778_),
    .B(_01785_),
    .X(_01786_));
 sky130_fd_sc_hd__mux2_1 _06695_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01787_));
 sky130_fd_sc_hd__o21a_1 _06696_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_01787_),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _06697_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _06698_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_01790_));
 sky130_fd_sc_hd__o21ba_1 _06699_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_01790_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(_01791_));
 sky130_fd_sc_hd__o21a_1 _06700_ (.A1(_01778_),
    .A2(_01789_),
    .B1(_01791_),
    .X(_01792_));
 sky130_fd_sc_hd__a211oi_1 _06701_ (.A1(_01786_),
    .A2(_01788_),
    .B1(_01792_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .Y(_01793_));
 sky130_fd_sc_hd__a31o_1 _06702_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .A2(_01780_),
    .A3(_01784_),
    .B1(_01793_),
    .X(_01794_));
 sky130_fd_sc_hd__and2b_1 _06703_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .X(_01795_));
 sky130_fd_sc_hd__a21bo_1 _06704_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01796_));
 sky130_fd_sc_hd__mux2_1 _06705_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .X(_01797_));
 sky130_fd_sc_hd__o221a_1 _06706_ (.A1(_01795_),
    .A2(_01796_),
    .B1(_01797_),
    .B2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .X(_01798_));
 sky130_fd_sc_hd__inv_2 _06707_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .Y(_01799_));
 sky130_fd_sc_hd__mux4_1 _06708_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01800_));
 sky130_fd_sc_hd__a21bo_1 _06709_ (.A1(_01799_),
    .A2(_01800_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .X(_01801_));
 sky130_fd_sc_hd__mux4_1 _06710_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01802_));
 sky130_fd_sc_hd__mux4_1 _06711_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _06712_ (.A0(_01802_),
    .A1(_01803_),
    .S(_01799_),
    .X(_01804_));
 sky130_fd_sc_hd__o22a_4 _06713_ (.A1(_01798_),
    .A2(_01801_),
    .B1(_01804_),
    .B2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _06714_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ),
    .S(_01805_),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _06715_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ),
    .S(_01805_),
    .X(_01807_));
 sky130_fd_sc_hd__mux4_1 _06716_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _06717_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(_01809_));
 sky130_fd_sc_hd__and2b_1 _06718_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .B(_01809_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _06719_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(_01811_));
 sky130_fd_sc_hd__a21bo_1 _06720_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .A2(_01811_),
    .B1_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(_01812_));
 sky130_fd_sc_hd__o221a_1 _06721_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .A2(_01808_),
    .B1(_01810_),
    .B2(_01812_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .X(_01813_));
 sky130_fd_sc_hd__mux4_1 _06722_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_01814_));
 sky130_fd_sc_hd__mux4_1 _06723_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _06724_ (.A0(_01814_),
    .A1(_01815_),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(_01816_));
 sky130_fd_sc_hd__and2b_1 _06725_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .B(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__nor2_2 _06726_ (.A(_01813_),
    .B(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__mux2_1 _06727_ (.A0(_01806_),
    .A1(_01807_),
    .S(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _06728_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ),
    .S(_01805_),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _06729_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ),
    .S(_01805_),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _06730_ (.A0(_01820_),
    .A1(_01821_),
    .S(_01818_),
    .X(_01822_));
 sky130_fd_sc_hd__inv_2 _06731_ (.A(net3845),
    .Y(_01823_));
 sky130_fd_sc_hd__mux4_1 _06732_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01824_));
 sky130_fd_sc_hd__mux4_1 _06733_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _06734_ (.A0(_01824_),
    .A1(_01825_),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .X(_01826_));
 sky130_fd_sc_hd__inv_2 _06735_ (.A(net3993),
    .Y(_01827_));
 sky130_fd_sc_hd__or2_1 _06736_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(_01828_));
 sky130_fd_sc_hd__o211a_1 _06737_ (.A1(_01827_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.half_q ),
    .B1(_01828_),
    .C1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01829_));
 sky130_fd_sc_hd__inv_2 _06738_ (.A(net3861),
    .Y(_01830_));
 sky130_fd_sc_hd__mux2_1 _06739_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(_01831_));
 sky130_fd_sc_hd__inv_2 _06740_ (.A(net3552),
    .Y(_01832_));
 sky130_fd_sc_hd__a21o_1 _06741_ (.A1(_01830_),
    .A2(_01831_),
    .B1(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__mux4_1 _06742_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_01834_));
 sky130_fd_sc_hd__or2_1 _06743_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .B(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__o211a_1 _06744_ (.A1(_01829_),
    .A2(_01833_),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ),
    .C1(_01835_),
    .X(_01836_));
 sky130_fd_sc_hd__a21oi_2 _06745_ (.A1(_01823_),
    .A2(_01826_),
    .B1(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__mux2_1 _06746_ (.A0(_01819_),
    .A1(_01822_),
    .S(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_1 _06747_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ),
    .S(_01805_),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _06748_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ),
    .S(_01805_),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _06749_ (.A0(_01839_),
    .A1(_01840_),
    .S(_01818_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _06750_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ),
    .S(_01805_),
    .X(_01842_));
 sky130_fd_sc_hd__or3_1 _06751_ (.A(_01813_),
    .B(_01817_),
    .C(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _06752_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ),
    .S(_01805_),
    .X(_01844_));
 sky130_fd_sc_hd__o21ba_1 _06753_ (.A1(_01818_),
    .A2(_01844_),
    .B1_N(_01837_),
    .X(_01845_));
 sky130_fd_sc_hd__a31oi_1 _06754_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .A2(_01780_),
    .A3(_01784_),
    .B1(_01793_),
    .Y(_01846_));
 sky130_fd_sc_hd__a221o_1 _06755_ (.A1(_01837_),
    .A2(_01841_),
    .B1(_01843_),
    .B2(_01845_),
    .C1(_01846_),
    .X(_01847_));
 sky130_fd_sc_hd__o211ai_4 _06756_ (.A1(_01794_),
    .A2(_01838_),
    .B1(_01847_),
    .C1(_01578_),
    .Y(_01848_));
 sky130_fd_sc_hd__a22o_4 _06757_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .A2(_01775_),
    .B1(_01776_),
    .B2(_01848_),
    .X(_01849_));
 sky130_fd_sc_hd__clkinv_2 _06758_ (.A(_01849_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__clkbuf_4 _06759_ (.A(_00188_),
    .X(_01850_));
 sky130_fd_sc_hd__buf_6 _06760_ (.A(_00220_),
    .X(_01851_));
 sky130_fd_sc_hd__a221o_1 _06761_ (.A1(_01850_),
    .A2(_01763_),
    .B1(_01765_),
    .B2(net3175),
    .C1(_01851_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__inv_2 _06762_ (.A(net3727),
    .Y(_01852_));
 sky130_fd_sc_hd__mux4_1 _06763_ (.A0(_01678_),
    .A1(_01585_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A3(_01676_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .S1(_01852_),
    .X(_01853_));
 sky130_fd_sc_hd__mux4_1 _06764_ (.A0(_01584_),
    .A1(_01587_),
    .A2(_01589_),
    .A3(_01590_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .S1(net4219),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _06765_ (.A0(_01853_),
    .A1(_01854_),
    .S(net3655),
    .X(_01855_));
 sky130_fd_sc_hd__clkbuf_1 _06766_ (.A(_01855_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ));
 sky130_fd_sc_hd__nor2_1 _06767_ (.A(_01332_),
    .B(_01388_),
    .Y(_01856_));
 sky130_fd_sc_hd__o221a_1 _06768_ (.A1(_01389_),
    .A2(_01390_),
    .B1(_01391_),
    .B2(_01356_),
    .C1(_01332_),
    .X(_01857_));
 sky130_fd_sc_hd__buf_8 _06769_ (.A(_01578_),
    .X(_01858_));
 sky130_fd_sc_hd__o21a_1 _06770_ (.A1(_01856_),
    .A2(_01857_),
    .B1(_01858_),
    .X(_01859_));
 sky130_fd_sc_hd__a22o_1 _06771_ (.A1(_00865_),
    .A2(_00869_),
    .B1(_00872_),
    .B2(_00811_),
    .X(_01860_));
 sky130_fd_sc_hd__and2_1 _06772_ (.A(_01858_),
    .B(_01860_),
    .X(_01861_));
 sky130_fd_sc_hd__nand2_2 _06773_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.m[0] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.m[1] ),
    .Y(_01862_));
 sky130_fd_sc_hd__buf_8 _06774_ (.A(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _06775_ (.A0(_01859_),
    .A1(_01861_),
    .S(_01863_),
    .X(_01864_));
 sky130_fd_sc_hd__clkbuf_1 _06776_ (.A(_01864_),
    .X(_00012_));
 sky130_fd_sc_hd__mux4_1 _06777_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A2(_01584_),
    .A3(_01585_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .X(_01865_));
 sky130_fd_sc_hd__mux4_1 _06778_ (.A0(_01587_),
    .A1(_01588_),
    .A2(_01589_),
    .A3(_01590_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _06779_ (.A0(_01865_),
    .A1(_01866_),
    .S(net3676),
    .X(_01867_));
 sky130_fd_sc_hd__clkbuf_1 _06780_ (.A(_01867_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ));
 sky130_fd_sc_hd__mux4_1 _06781_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(_01676_),
    .A2(_01587_),
    .A3(_01588_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(_01868_));
 sky130_fd_sc_hd__mux4_1 _06782_ (.A0(_01678_),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(_01589_),
    .A3(_01590_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _06783_ (.A0(_01868_),
    .A1(_01869_),
    .S(net3262),
    .X(_01870_));
 sky130_fd_sc_hd__clkbuf_1 _06784_ (.A(net3263),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ));
 sky130_fd_sc_hd__mux4_1 _06785_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A1(_01676_),
    .A2(_01678_),
    .A3(_01585_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .X(_01871_));
 sky130_fd_sc_hd__mux4_1 _06786_ (.A0(_01584_),
    .A1(_01588_),
    .A2(_01589_),
    .A3(_01590_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .X(_01872_));
 sky130_fd_sc_hd__mux2_1 _06787_ (.A0(_01871_),
    .A1(_01872_),
    .S(net3654),
    .X(_01873_));
 sky130_fd_sc_hd__clkbuf_1 _06788_ (.A(_01873_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ));
 sky130_fd_sc_hd__mux4_1 _06789_ (.A0(_01584_),
    .A1(_01587_),
    .A2(_01589_),
    .A3(_01590_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .X(_01874_));
 sky130_fd_sc_hd__mux4_1 _06790_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A3(_01585_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .X(_01875_));
 sky130_fd_sc_hd__inv_2 _06791_ (.A(net3404),
    .Y(_01876_));
 sky130_fd_sc_hd__mux2_1 _06792_ (.A0(_01874_),
    .A1(_01875_),
    .S(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__clkbuf_1 _06793_ (.A(net3405),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ));
 sky130_fd_sc_hd__buf_8 _06794_ (.A(_00311_),
    .X(_01878_));
 sky130_fd_sc_hd__nand3b_2 _06795_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .C(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__or3_1 _06796_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_01880_));
 sky130_fd_sc_hd__or2_1 _06797_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__clkbuf_2 _06798_ (.A(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__o21a_2 _06799_ (.A1(_01879_),
    .A2(_01882_),
    .B1(_00408_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _06800_ (.A0(_01495_),
    .A1(net3293),
    .S(_01883_),
    .X(_01884_));
 sky130_fd_sc_hd__clkbuf_1 _06801_ (.A(_01884_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _06802_ (.A0(_01500_),
    .A1(net3588),
    .S(_01883_),
    .X(_01885_));
 sky130_fd_sc_hd__clkbuf_1 _06803_ (.A(_01885_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _06804_ (.A0(_01581_),
    .A1(net3478),
    .S(_01883_),
    .X(_01886_));
 sky130_fd_sc_hd__clkbuf_1 _06805_ (.A(_01886_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _06806_ (.A0(_01423_),
    .A1(net3528),
    .S(_01883_),
    .X(_01887_));
 sky130_fd_sc_hd__clkbuf_1 _06807_ (.A(_01887_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _06808_ (.A(net4147),
    .X(_01888_));
 sky130_fd_sc_hd__clkbuf_2 _06809_ (.A(net4149),
    .X(_01889_));
 sky130_fd_sc_hd__inv_2 _06810_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .Y(_01890_));
 sky130_fd_sc_hd__or4_1 _06811_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_01889_),
    .C(_01890_),
    .D(_01879_),
    .X(_01891_));
 sky130_fd_sc_hd__o21a_2 _06812_ (.A1(_01888_),
    .A2(_01891_),
    .B1(_00408_),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _06813_ (.A0(_01495_),
    .A1(net3696),
    .S(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__clkbuf_1 _06814_ (.A(_01893_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _06815_ (.A0(_01500_),
    .A1(net3453),
    .S(_01892_),
    .X(_01894_));
 sky130_fd_sc_hd__clkbuf_1 _06816_ (.A(_01894_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _06817_ (.A0(_01581_),
    .A1(net3301),
    .S(_01892_),
    .X(_01895_));
 sky130_fd_sc_hd__clkbuf_1 _06818_ (.A(_01895_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _06819_ (.A0(_01423_),
    .A1(net3319),
    .S(_01892_),
    .X(_01896_));
 sky130_fd_sc_hd__clkbuf_1 _06820_ (.A(_01896_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__clkinv_2 _06821_ (.A(net3601),
    .Y(_01897_));
 sky130_fd_sc_hd__nand2_1 _06822_ (.A(_00171_),
    .B(_01882_),
    .Y(_01898_));
 sky130_fd_sc_hd__inv_2 _06823_ (.A(_01888_),
    .Y(_01899_));
 sky130_fd_sc_hd__or3_1 _06824_ (.A(_01889_),
    .B(_01899_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_01900_));
 sky130_fd_sc_hd__inv_2 _06825_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .Y(_01901_));
 sky130_fd_sc_hd__and3b_1 _06826_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .C(_01415_),
    .X(_01902_));
 sky130_fd_sc_hd__and3b_1 _06827_ (.A_N(_01900_),
    .B(_01901_),
    .C(_01902_),
    .X(_01903_));
 sky130_fd_sc_hd__mux2_1 _06828_ (.A0(_01897_),
    .A1(_01898_),
    .S(_01903_),
    .X(_01904_));
 sky130_fd_sc_hd__o21ai_1 _06829_ (.A1(_00646_),
    .A2(_01904_),
    .B1(_00614_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__buf_2 _06830_ (.A(_00363_),
    .X(_01905_));
 sky130_fd_sc_hd__inv_2 _06831_ (.A(net3557),
    .Y(_01906_));
 sky130_fd_sc_hd__nand2_1 _06832_ (.A(_01446_),
    .B(_01882_),
    .Y(_01907_));
 sky130_fd_sc_hd__mux2_1 _06833_ (.A0(_01906_),
    .A1(_01907_),
    .S(_01903_),
    .X(_01908_));
 sky130_fd_sc_hd__o21ai_1 _06834_ (.A1(_01905_),
    .A2(_01908_),
    .B1(_01481_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__inv_2 _06835_ (.A(net3398),
    .Y(_01909_));
 sky130_fd_sc_hd__nand2_1 _06836_ (.A(_00551_),
    .B(_01882_),
    .Y(_01910_));
 sky130_fd_sc_hd__mux2_1 _06837_ (.A0(_01909_),
    .A1(_01910_),
    .S(_01903_),
    .X(_01911_));
 sky130_fd_sc_hd__buf_4 _06838_ (.A(_00251_),
    .X(_01912_));
 sky130_fd_sc_hd__o21ai_1 _06839_ (.A1(_01905_),
    .A2(_01911_),
    .B1(_01912_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__inv_2 _06840_ (.A(net3407),
    .Y(_01913_));
 sky130_fd_sc_hd__nand2_2 _06841_ (.A(_01452_),
    .B(_01882_),
    .Y(_01914_));
 sky130_fd_sc_hd__mux2_1 _06842_ (.A0(_01913_),
    .A1(_01914_),
    .S(_01903_),
    .X(_01915_));
 sky130_fd_sc_hd__o21ai_1 _06843_ (.A1(_01905_),
    .A2(_01915_),
    .B1(_00621_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _06844_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_01879_),
    .Y(_01916_));
 sky130_fd_sc_hd__and3b_1 _06845_ (.A_N(_01889_),
    .B(_01888_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_01917_));
 sky130_fd_sc_hd__a21oi_4 _06846_ (.A1(_01916_),
    .A2(_01917_),
    .B1(_00267_),
    .Y(_01918_));
 sky130_fd_sc_hd__mux2_1 _06847_ (.A0(_01495_),
    .A1(net3336),
    .S(_01918_),
    .X(_01919_));
 sky130_fd_sc_hd__clkbuf_1 _06848_ (.A(_01919_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _06849_ (.A0(_01500_),
    .A1(net3519),
    .S(_01918_),
    .X(_01920_));
 sky130_fd_sc_hd__clkbuf_1 _06850_ (.A(_01920_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _06851_ (.A0(_01581_),
    .A1(net3526),
    .S(_01918_),
    .X(_01921_));
 sky130_fd_sc_hd__clkbuf_1 _06852_ (.A(_01921_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _06853_ (.A0(_01423_),
    .A1(net3662),
    .S(_01918_),
    .X(_01922_));
 sky130_fd_sc_hd__clkbuf_1 _06854_ (.A(_01922_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__clkbuf_4 _06855_ (.A(_00196_),
    .X(_01923_));
 sky130_fd_sc_hd__and4_1 _06856_ (.A(_01889_),
    .B(_01899_),
    .C(_01890_),
    .D(_01916_),
    .X(_01924_));
 sky130_fd_sc_hd__clkbuf_2 _06857_ (.A(_01924_),
    .X(_01925_));
 sky130_fd_sc_hd__or2_1 _06858_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .B(_01925_),
    .X(_01926_));
 sky130_fd_sc_hd__nand2_1 _06859_ (.A(_01898_),
    .B(_01925_),
    .Y(_01927_));
 sky130_fd_sc_hd__a31o_1 _06860_ (.A1(_01923_),
    .A2(_01926_),
    .A3(_01927_),
    .B1(_00603_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__or2_1 _06861_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .B(_01925_),
    .X(_01928_));
 sky130_fd_sc_hd__nand2_1 _06862_ (.A(_01907_),
    .B(_01925_),
    .Y(_01929_));
 sky130_fd_sc_hd__a31o_1 _06863_ (.A1(_01923_),
    .A2(_01928_),
    .A3(_01929_),
    .B1(_00487_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__or2_1 _06864_ (.A(net4142),
    .B(_01925_),
    .X(_01930_));
 sky130_fd_sc_hd__nand2_1 _06865_ (.A(_01910_),
    .B(_01925_),
    .Y(_01931_));
 sky130_fd_sc_hd__a31o_1 _06866_ (.A1(_01923_),
    .A2(_01930_),
    .A3(_01931_),
    .B1(_00394_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _06867_ (.A(net4089),
    .B(_01925_),
    .Y(_01932_));
 sky130_fd_sc_hd__a211o_1 _06868_ (.A1(_01914_),
    .A2(_01925_),
    .B1(_01932_),
    .C1(_01471_),
    .X(_01933_));
 sky130_fd_sc_hd__nand2_1 _06869_ (.A(_00263_),
    .B(_01933_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _06870_ (.A1(_01889_),
    .A2(_01899_),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .A4(_01916_),
    .B1(_00522_),
    .X(_01934_));
 sky130_fd_sc_hd__mux2_1 _06871_ (.A0(net4110),
    .A1(_00692_),
    .S(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__clkbuf_1 _06872_ (.A(_01935_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _06873_ (.A0(net4032),
    .A1(_00695_),
    .S(_01934_),
    .X(_01936_));
 sky130_fd_sc_hd__clkbuf_1 _06874_ (.A(_01936_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _06875_ (.A0(net3980),
    .A1(_00697_),
    .S(_01934_),
    .X(_01937_));
 sky130_fd_sc_hd__clkbuf_1 _06876_ (.A(_01937_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _06877_ (.A0(net3692),
    .A1(_00528_),
    .S(_01934_),
    .X(_01938_));
 sky130_fd_sc_hd__clkbuf_1 _06878_ (.A(_01938_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_1 _06879_ (.A(_01889_),
    .B(_01888_),
    .C(_01890_),
    .D(_01916_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _06880_ (.A0(_00948_),
    .A1(_01898_),
    .S(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__o21ai_1 _06881_ (.A1(_01905_),
    .A2(_01940_),
    .B1(_00614_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _06882_ (.A0(_00951_),
    .A1(_01907_),
    .S(_01939_),
    .X(_01941_));
 sky130_fd_sc_hd__o21ai_1 _06883_ (.A1(_01905_),
    .A2(_01941_),
    .B1(_01481_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _06884_ (.A0(_00953_),
    .A1(_01910_),
    .S(_01939_),
    .X(_01942_));
 sky130_fd_sc_hd__o21ai_1 _06885_ (.A1(_01905_),
    .A2(_01942_),
    .B1(_01912_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _06886_ (.A0(_00943_),
    .A1(_01914_),
    .S(_01939_),
    .X(_01943_));
 sky130_fd_sc_hd__o21ai_1 _06887_ (.A1(_01905_),
    .A2(_01943_),
    .B1(_00621_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _06888_ (.A1(_01889_),
    .A2(_01888_),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .A4(_01916_),
    .B1(_00522_),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_1 _06889_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .A1(_00692_),
    .S(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__clkbuf_1 _06890_ (.A(_01945_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _06891_ (.A0(net3960),
    .A1(_00695_),
    .S(_01944_),
    .X(_01946_));
 sky130_fd_sc_hd__clkbuf_1 _06892_ (.A(_01946_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _06893_ (.A0(net3644),
    .A1(_00697_),
    .S(_01944_),
    .X(_01947_));
 sky130_fd_sc_hd__clkbuf_1 _06894_ (.A(_01947_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _06895_ (.A0(net4071),
    .A1(_00528_),
    .S(_01944_),
    .X(_01948_));
 sky130_fd_sc_hd__clkbuf_1 _06896_ (.A(_01948_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__o31a_2 _06897_ (.A1(_01901_),
    .A2(_01879_),
    .A3(_01880_),
    .B1(_01489_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _06898_ (.A0(_01495_),
    .A1(net3919),
    .S(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__clkbuf_1 _06899_ (.A(_01950_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _06900_ (.A0(_01500_),
    .A1(net3195),
    .S(_01949_),
    .X(_01951_));
 sky130_fd_sc_hd__clkbuf_1 _06901_ (.A(_01951_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _06902_ (.A0(_01581_),
    .A1(net3581),
    .S(_01949_),
    .X(_01952_));
 sky130_fd_sc_hd__clkbuf_1 _06903_ (.A(_01952_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _06904_ (.A0(_01423_),
    .A1(net3372),
    .S(_01949_),
    .X(_01953_));
 sky130_fd_sc_hd__clkbuf_1 _06905_ (.A(_01953_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__nand2_1 _06906_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_01880_),
    .Y(_01954_));
 sky130_fd_sc_hd__a21o_1 _06907_ (.A1(_01882_),
    .A2(_01954_),
    .B1(_01879_),
    .X(_01955_));
 sky130_fd_sc_hd__o41a_2 _06908_ (.A1(_01889_),
    .A2(_01888_),
    .A3(_01890_),
    .A4(_01955_),
    .B1(_01497_),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_1 _06909_ (.A0(_01495_),
    .A1(net3918),
    .S(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__clkbuf_1 _06910_ (.A(_01957_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _06911_ (.A0(_01500_),
    .A1(net3321),
    .S(_01956_),
    .X(_01958_));
 sky130_fd_sc_hd__clkbuf_1 _06912_ (.A(_01958_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _06913_ (.A0(_01581_),
    .A1(net3990),
    .S(_01956_),
    .X(_01959_));
 sky130_fd_sc_hd__clkbuf_1 _06914_ (.A(_01959_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _06915_ (.A0(_01423_),
    .A1(net3682),
    .S(_01956_),
    .X(_01960_));
 sky130_fd_sc_hd__clkbuf_1 _06916_ (.A(_01960_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__inv_2 _06917_ (.A(net3595),
    .Y(_01961_));
 sky130_fd_sc_hd__nor2_2 _06918_ (.A(_01900_),
    .B(_01955_),
    .Y(_01962_));
 sky130_fd_sc_hd__mux2_1 _06919_ (.A0(_01961_),
    .A1(_01898_),
    .S(_01962_),
    .X(_01963_));
 sky130_fd_sc_hd__o21ai_1 _06920_ (.A1(_01905_),
    .A2(_01963_),
    .B1(_00614_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__nand2_1 _06921_ (.A(_01907_),
    .B(_01962_),
    .Y(_01964_));
 sky130_fd_sc_hd__or2_1 _06922_ (.A(net4191),
    .B(_01962_),
    .X(_01965_));
 sky130_fd_sc_hd__a31o_1 _06923_ (.A1(_01923_),
    .A2(_01964_),
    .A3(_01965_),
    .B1(_00487_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__inv_2 _06924_ (.A(net3628),
    .Y(_01966_));
 sky130_fd_sc_hd__mux2_1 _06925_ (.A0(_01966_),
    .A1(_01910_),
    .S(_01962_),
    .X(_01967_));
 sky130_fd_sc_hd__o21ai_1 _06926_ (.A1(_01905_),
    .A2(_01967_),
    .B1(_01912_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__inv_2 _06927_ (.A(net3802),
    .Y(_01968_));
 sky130_fd_sc_hd__mux2_1 _06928_ (.A0(_01968_),
    .A1(_01914_),
    .S(_01962_),
    .X(_01969_));
 sky130_fd_sc_hd__o21ai_1 _06929_ (.A1(_01905_),
    .A2(_01969_),
    .B1(_00621_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3_2 _06930_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_01902_),
    .C(_01917_),
    .X(_01970_));
 sky130_fd_sc_hd__clkbuf_4 _06931_ (.A(_00181_),
    .X(_01971_));
 sky130_fd_sc_hd__nor2_1 _06932_ (.A(_01971_),
    .B(_01970_),
    .Y(_01972_));
 sky130_fd_sc_hd__a221o_1 _06933_ (.A1(_01762_),
    .A2(_01970_),
    .B1(_01972_),
    .B2(net3340),
    .C1(_01766_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _06934_ (.A1(_01771_),
    .A2(_01970_),
    .B1(_01972_),
    .B2(net3230),
    .C1(_01772_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__clkbuf_4 _06935_ (.A(_00221_),
    .X(_01973_));
 sky130_fd_sc_hd__a221o_1 _06936_ (.A1(_01850_),
    .A2(_01970_),
    .B1(_01972_),
    .B2(net3194),
    .C1(_01973_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__a22o_1 _06937_ (.A1(_00960_),
    .A2(_00962_),
    .B1(_00965_),
    .B2(_00956_),
    .X(_01974_));
 sky130_fd_sc_hd__and2_1 _06938_ (.A(_01858_),
    .B(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_1 _06939_ (.A0(_01861_),
    .A1(_01975_),
    .S(_01863_),
    .X(_01976_));
 sky130_fd_sc_hd__clkbuf_1 _06940_ (.A(_01976_),
    .X(_00013_));
 sky130_fd_sc_hd__nand3b_2 _06941_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .C(_01878_),
    .Y(_01977_));
 sky130_fd_sc_hd__or3_1 _06942_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_01978_));
 sky130_fd_sc_hd__or2_2 _06943_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__o21a_2 _06944_ (.A1(_01977_),
    .A2(_01979_),
    .B1(_00408_),
    .X(_01980_));
 sky130_fd_sc_hd__mux2_1 _06945_ (.A0(_01495_),
    .A1(net3411),
    .S(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__clkbuf_1 _06946_ (.A(_01981_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _06947_ (.A0(_01500_),
    .A1(net3315),
    .S(_01980_),
    .X(_01982_));
 sky130_fd_sc_hd__clkbuf_1 _06948_ (.A(_01982_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _06949_ (.A0(_01581_),
    .A1(net3748),
    .S(_01980_),
    .X(_01983_));
 sky130_fd_sc_hd__clkbuf_1 _06950_ (.A(_01983_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__buf_4 _06951_ (.A(_00191_),
    .X(_01984_));
 sky130_fd_sc_hd__mux2_1 _06952_ (.A0(_01984_),
    .A1(net3587),
    .S(_01980_),
    .X(_01985_));
 sky130_fd_sc_hd__clkbuf_1 _06953_ (.A(_01985_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__inv_2 _06954_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .Y(_01986_));
 sky130_fd_sc_hd__and3b_1 _06955_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .C(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ),
    .X(_01987_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06956_ (.A(_01987_),
    .X(_01988_));
 sky130_fd_sc_hd__nand2_1 _06957_ (.A(_01986_),
    .B(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__clkbuf_2 _06958_ (.A(net4140),
    .X(_01990_));
 sky130_fd_sc_hd__or3b_1 _06959_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(_01990_),
    .C_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_01991_));
 sky130_fd_sc_hd__o21a_2 _06960_ (.A1(_01989_),
    .A2(_01991_),
    .B1(_00408_),
    .X(_01992_));
 sky130_fd_sc_hd__mux2_1 _06961_ (.A0(_01495_),
    .A1(net3428),
    .S(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__clkbuf_1 _06962_ (.A(_01993_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _06963_ (.A0(_01500_),
    .A1(net3510),
    .S(_01992_),
    .X(_01994_));
 sky130_fd_sc_hd__clkbuf_1 _06964_ (.A(_01994_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _06965_ (.A0(_01581_),
    .A1(net3604),
    .S(_01992_),
    .X(_01995_));
 sky130_fd_sc_hd__clkbuf_1 _06966_ (.A(_01995_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _06967_ (.A0(_01984_),
    .A1(net3704),
    .S(_01992_),
    .X(_01996_));
 sky130_fd_sc_hd__clkbuf_1 _06968_ (.A(_01996_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__clkbuf_4 _06969_ (.A(_00363_),
    .X(_01997_));
 sky130_fd_sc_hd__inv_2 _06970_ (.A(_01990_),
    .Y(_01998_));
 sky130_fd_sc_hd__or3_2 _06971_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(_01998_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_01999_));
 sky130_fd_sc_hd__nand2_1 _06972_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_01978_),
    .Y(_02000_));
 sky130_fd_sc_hd__and2_1 _06973_ (.A(_01979_),
    .B(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__nand2_1 _06974_ (.A(_01988_),
    .B(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hd__buf_8 _06975_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[0] ),
    .X(_02003_));
 sky130_fd_sc_hd__nand2_1 _06976_ (.A(_02003_),
    .B(_01979_),
    .Y(_02004_));
 sky130_fd_sc_hd__or2_1 _06977_ (.A(_01989_),
    .B(_01999_),
    .X(_02005_));
 sky130_fd_sc_hd__nand2_1 _06978_ (.A(net3540),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__o31a_1 _06979_ (.A1(_01999_),
    .A2(_02002_),
    .A3(_02004_),
    .B1(_02006_),
    .X(_02007_));
 sky130_fd_sc_hd__o21ai_1 _06980_ (.A1(_01997_),
    .A2(_02007_),
    .B1(_00614_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_1 _06981_ (.A(_01446_),
    .B(_01979_),
    .Y(_02008_));
 sky130_fd_sc_hd__nand2_1 _06982_ (.A(net3570),
    .B(_02005_),
    .Y(_02009_));
 sky130_fd_sc_hd__o31a_1 _06983_ (.A1(_01999_),
    .A2(_02002_),
    .A3(_02008_),
    .B1(_02009_),
    .X(_02010_));
 sky130_fd_sc_hd__o21ai_1 _06984_ (.A1(_01997_),
    .A2(_02010_),
    .B1(_01481_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__and2_1 _06985_ (.A(_00187_),
    .B(_01979_),
    .X(_02011_));
 sky130_fd_sc_hd__nor2_1 _06986_ (.A(_01989_),
    .B(_01999_),
    .Y(_02012_));
 sky130_fd_sc_hd__mux2_1 _06987_ (.A0(net3686),
    .A1(_02011_),
    .S(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__a21o_1 _06988_ (.A1(_00279_),
    .A2(_02013_),
    .B1(_00222_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__inv_2 _06989_ (.A(net3640),
    .Y(_02014_));
 sky130_fd_sc_hd__nand2_1 _06990_ (.A(_01452_),
    .B(_01979_),
    .Y(_02015_));
 sky130_fd_sc_hd__mux2_1 _06991_ (.A0(_02014_),
    .A1(_02015_),
    .S(_02012_),
    .X(_02016_));
 sky130_fd_sc_hd__o21ai_1 _06992_ (.A1(_01997_),
    .A2(_02016_),
    .B1(_00621_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _06993_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_01977_),
    .Y(_02017_));
 sky130_fd_sc_hd__and3b_1 _06994_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(_01990_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_02018_));
 sky130_fd_sc_hd__a21oi_4 _06995_ (.A1(_02017_),
    .A2(_02018_),
    .B1(_00267_),
    .Y(_02019_));
 sky130_fd_sc_hd__mux2_1 _06996_ (.A0(_01495_),
    .A1(net3472),
    .S(_02019_),
    .X(_02020_));
 sky130_fd_sc_hd__clkbuf_1 _06997_ (.A(_02020_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _06998_ (.A0(_01500_),
    .A1(net3224),
    .S(_02019_),
    .X(_02021_));
 sky130_fd_sc_hd__clkbuf_1 _06999_ (.A(_02021_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _07000_ (.A0(_01581_),
    .A1(net3530),
    .S(_02019_),
    .X(_02022_));
 sky130_fd_sc_hd__clkbuf_1 _07001_ (.A(_02022_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _07002_ (.A0(_01984_),
    .A1(net3274),
    .S(_02019_),
    .X(_02023_));
 sky130_fd_sc_hd__clkbuf_1 _07003_ (.A(_02023_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4bb_2 _07004_ (.A_N(_01990_),
    .B_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .C(_02017_),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .X(_02024_));
 sky130_fd_sc_hd__nand2_1 _07005_ (.A(_02004_),
    .B(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__or2_1 _07006_ (.A(net4195),
    .B(_02024_),
    .X(_02026_));
 sky130_fd_sc_hd__a31o_1 _07007_ (.A1(_01923_),
    .A2(_02025_),
    .A3(_02026_),
    .B1(_00603_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _07008_ (.A(_02008_),
    .B(_02024_),
    .Y(_02027_));
 sky130_fd_sc_hd__or2_1 _07009_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .B(_02024_),
    .X(_02028_));
 sky130_fd_sc_hd__a31o_1 _07010_ (.A1(_01923_),
    .A2(_02027_),
    .A3(_02028_),
    .B1(_00487_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__or2b_1 _07011_ (.A(_02011_),
    .B_N(_02024_),
    .X(_02029_));
 sky130_fd_sc_hd__or2_1 _07012_ (.A(net4143),
    .B(_02024_),
    .X(_02030_));
 sky130_fd_sc_hd__a31o_1 _07013_ (.A1(_01923_),
    .A2(_02029_),
    .A3(_02030_),
    .B1(_00394_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__buf_6 _07014_ (.A(_00227_),
    .X(_02031_));
 sky130_fd_sc_hd__nor2_1 _07015_ (.A(net3985),
    .B(_02024_),
    .Y(_02032_));
 sky130_fd_sc_hd__a211o_1 _07016_ (.A1(_02015_),
    .A2(_02024_),
    .B1(_02032_),
    .C1(_01471_),
    .X(_02033_));
 sky130_fd_sc_hd__nand2_1 _07017_ (.A(_02031_),
    .B(_02033_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__clkbuf_4 _07018_ (.A(_00180_),
    .X(_02034_));
 sky130_fd_sc_hd__a41o_2 _07019_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .A2(_01998_),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .A4(_02017_),
    .B1(_02034_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _07020_ (.A0(net4067),
    .A1(_00692_),
    .S(_02035_),
    .X(_02036_));
 sky130_fd_sc_hd__clkbuf_1 _07021_ (.A(_02036_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _07022_ (.A0(net4210),
    .A1(_00695_),
    .S(_02035_),
    .X(_02037_));
 sky130_fd_sc_hd__clkbuf_1 _07023_ (.A(_02037_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _07024_ (.A0(net4014),
    .A1(_00697_),
    .S(_02035_),
    .X(_02038_));
 sky130_fd_sc_hd__clkbuf_1 _07025_ (.A(_02038_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _07026_ (.A0(net3873),
    .A1(_00528_),
    .S(_02035_),
    .X(_02039_));
 sky130_fd_sc_hd__clkbuf_1 _07027_ (.A(_02039_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4b_2 _07028_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .B(_02017_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .D(_01990_),
    .X(_02040_));
 sky130_fd_sc_hd__or2_1 _07029_ (.A(net4206),
    .B(_02040_),
    .X(_02041_));
 sky130_fd_sc_hd__nand2_1 _07030_ (.A(_02004_),
    .B(_02040_),
    .Y(_02042_));
 sky130_fd_sc_hd__a31o_1 _07031_ (.A1(_01923_),
    .A2(_02041_),
    .A3(_02042_),
    .B1(_00603_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _07032_ (.A0(_01246_),
    .A1(_02008_),
    .S(_02040_),
    .X(_02043_));
 sky130_fd_sc_hd__o21ai_1 _07033_ (.A1(_01997_),
    .A2(_02043_),
    .B1(_01481_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__buf_6 _07034_ (.A(_00196_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _07035_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .A1(_02011_),
    .S(_02040_),
    .X(_02045_));
 sky130_fd_sc_hd__a21o_1 _07036_ (.A1(_02044_),
    .A2(_02045_),
    .B1(_00222_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _07037_ (.A0(_01238_),
    .A1(_02015_),
    .S(_02040_),
    .X(_02046_));
 sky130_fd_sc_hd__o21ai_1 _07038_ (.A1(_01997_),
    .A2(_02046_),
    .B1(_00621_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _07039_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .A2(_01990_),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .A4(_02017_),
    .B1(_02034_),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _07040_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .A1(_00692_),
    .S(_02047_),
    .X(_02048_));
 sky130_fd_sc_hd__clkbuf_1 _07041_ (.A(_02048_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _07042_ (.A0(net4041),
    .A1(_00695_),
    .S(_02047_),
    .X(_02049_));
 sky130_fd_sc_hd__clkbuf_1 _07043_ (.A(_02049_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _07044_ (.A0(net3502),
    .A1(_00697_),
    .S(_02047_),
    .X(_02050_));
 sky130_fd_sc_hd__clkbuf_1 _07045_ (.A(_02050_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__buf_6 _07046_ (.A(_00527_),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _07047_ (.A0(net4164),
    .A1(_02051_),
    .S(_02047_),
    .X(_02052_));
 sky130_fd_sc_hd__clkbuf_1 _07048_ (.A(_02052_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__o31a_2 _07049_ (.A1(_01986_),
    .A2(_01977_),
    .A3(_01978_),
    .B1(_01489_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _07050_ (.A0(_01495_),
    .A1(net3963),
    .S(_02053_),
    .X(_02054_));
 sky130_fd_sc_hd__clkbuf_1 _07051_ (.A(_02054_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _07052_ (.A0(_01500_),
    .A1(net3706),
    .S(_02053_),
    .X(_02055_));
 sky130_fd_sc_hd__clkbuf_1 _07053_ (.A(_02055_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _07054_ (.A0(_01581_),
    .A1(net3870),
    .S(_02053_),
    .X(_02056_));
 sky130_fd_sc_hd__clkbuf_1 _07055_ (.A(_02056_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _07056_ (.A0(_01984_),
    .A1(net3927),
    .S(_02053_),
    .X(_02057_));
 sky130_fd_sc_hd__clkbuf_1 _07057_ (.A(_02057_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__clkbuf_4 _07058_ (.A(_00171_),
    .X(_02058_));
 sky130_fd_sc_hd__or2_1 _07059_ (.A(_01977_),
    .B(_02001_),
    .X(_02059_));
 sky130_fd_sc_hd__o21a_1 _07060_ (.A1(_01991_),
    .A2(_02059_),
    .B1(_00408_),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _07061_ (.A0(_02058_),
    .A1(net3680),
    .S(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__clkbuf_1 _07062_ (.A(_02061_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__clkbuf_4 _07063_ (.A(_00184_),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_1 _07064_ (.A0(_02062_),
    .A1(net3515),
    .S(_02060_),
    .X(_02063_));
 sky130_fd_sc_hd__clkbuf_1 _07065_ (.A(_02063_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__clkbuf_4 _07066_ (.A(_00551_),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _07067_ (.A0(_02064_),
    .A1(net3759),
    .S(_02060_),
    .X(_02065_));
 sky130_fd_sc_hd__clkbuf_1 _07068_ (.A(_02065_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _07069_ (.A0(_01984_),
    .A1(net3285),
    .S(_02060_),
    .X(_02066_));
 sky130_fd_sc_hd__clkbuf_1 _07070_ (.A(_02066_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _07071_ (.A(_01999_),
    .B(_02059_),
    .Y(_02067_));
 sky130_fd_sc_hd__or2_1 _07072_ (.A(net3940),
    .B(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__nand2_1 _07073_ (.A(_02004_),
    .B(_02067_),
    .Y(_02069_));
 sky130_fd_sc_hd__a31o_1 _07074_ (.A1(_01923_),
    .A2(_02068_),
    .A3(_02069_),
    .B1(_00603_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__or2_1 _07075_ (.A(net4052),
    .B(_02067_),
    .X(_02070_));
 sky130_fd_sc_hd__nand2_1 _07076_ (.A(_02008_),
    .B(_02067_),
    .Y(_02071_));
 sky130_fd_sc_hd__a31o_1 _07077_ (.A1(_01923_),
    .A2(_02070_),
    .A3(_02071_),
    .B1(_00487_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__mux2_1 _07078_ (.A0(net3384),
    .A1(_02011_),
    .S(_02067_),
    .X(_02072_));
 sky130_fd_sc_hd__a21o_1 _07079_ (.A1(_02044_),
    .A2(_02072_),
    .B1(_00262_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__nor2_1 _07080_ (.A(net3849),
    .B(_02067_),
    .Y(_02073_));
 sky130_fd_sc_hd__a211o_1 _07081_ (.A1(_02015_),
    .A2(_02067_),
    .B1(_02073_),
    .C1(_01471_),
    .X(_02074_));
 sky130_fd_sc_hd__nand2_1 _07082_ (.A(_02031_),
    .B(_02074_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3_2 _07083_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_01988_),
    .C(_02018_),
    .X(_02075_));
 sky130_fd_sc_hd__nor2_1 _07084_ (.A(_01971_),
    .B(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__a221o_1 _07085_ (.A1(_01762_),
    .A2(_02075_),
    .B1(_02076_),
    .B2(net3289),
    .C1(_01766_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _07086_ (.A1(_01771_),
    .A2(_02075_),
    .B1(_02076_),
    .B2(net3187),
    .C1(_01772_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _07087_ (.A1(_01850_),
    .A2(_02075_),
    .B1(_02076_),
    .B2(net3259),
    .C1(_01973_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__and2_1 _07088_ (.A(_01858_),
    .B(_01309_),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_1 _07089_ (.A0(_01975_),
    .A1(_02077_),
    .S(_01863_),
    .X(_02078_));
 sky130_fd_sc_hd__clkbuf_1 _07090_ (.A(_02078_),
    .X(_00014_));
 sky130_fd_sc_hd__nand3b_2 _07091_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .C(_01878_),
    .Y(_02079_));
 sky130_fd_sc_hd__or3_1 _07092_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_02080_));
 sky130_fd_sc_hd__or2_1 _07093_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07094_ (.A(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__o21a_2 _07095_ (.A1(_02079_),
    .A2(_02082_),
    .B1(_00408_),
    .X(_02083_));
 sky130_fd_sc_hd__mux2_1 _07096_ (.A0(_02058_),
    .A1(net3805),
    .S(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__clkbuf_1 _07097_ (.A(_02084_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _07098_ (.A0(_02062_),
    .A1(net3771),
    .S(_02083_),
    .X(_02085_));
 sky130_fd_sc_hd__clkbuf_1 _07099_ (.A(_02085_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _07100_ (.A0(_02064_),
    .A1(net3750),
    .S(_02083_),
    .X(_02086_));
 sky130_fd_sc_hd__clkbuf_1 _07101_ (.A(_02086_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _07102_ (.A0(_01984_),
    .A1(net3823),
    .S(_02083_),
    .X(_02087_));
 sky130_fd_sc_hd__clkbuf_1 _07103_ (.A(_02087_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _07104_ (.A(net4170),
    .X(_02088_));
 sky130_fd_sc_hd__clkbuf_2 _07105_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .X(_02089_));
 sky130_fd_sc_hd__inv_2 _07106_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .Y(_02090_));
 sky130_fd_sc_hd__or4_1 _07107_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02089_),
    .C(_02090_),
    .D(_02079_),
    .X(_02091_));
 sky130_fd_sc_hd__buf_6 _07108_ (.A(_00407_),
    .X(_02092_));
 sky130_fd_sc_hd__o21a_2 _07109_ (.A1(_02088_),
    .A2(_02091_),
    .B1(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__mux2_1 _07110_ (.A0(_02058_),
    .A1(net3425),
    .S(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__clkbuf_1 _07111_ (.A(_02094_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _07112_ (.A0(_02062_),
    .A1(net3464),
    .S(_02093_),
    .X(_02095_));
 sky130_fd_sc_hd__clkbuf_1 _07113_ (.A(_02095_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _07114_ (.A0(_02064_),
    .A1(net3432),
    .S(_02093_),
    .X(_02096_));
 sky130_fd_sc_hd__clkbuf_1 _07115_ (.A(_02096_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _07116_ (.A0(_01984_),
    .A1(net3609),
    .S(_02093_),
    .X(_02097_));
 sky130_fd_sc_hd__clkbuf_1 _07117_ (.A(_02097_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _07118_ (.A(_02088_),
    .Y(_02098_));
 sky130_fd_sc_hd__or3_2 _07119_ (.A(_02089_),
    .B(_02098_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_02099_));
 sky130_fd_sc_hd__and3b_1 _07120_ (.A_N(\c.genblk1.genblk1.subs.cs[3].c.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .C(_00311_),
    .X(_02100_));
 sky130_fd_sc_hd__clkbuf_2 _07121_ (.A(_02100_),
    .X(_02101_));
 sky130_fd_sc_hd__nand2_1 _07122_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02080_),
    .Y(_02102_));
 sky130_fd_sc_hd__and2_1 _07123_ (.A(_02082_),
    .B(_02102_),
    .X(_02103_));
 sky130_fd_sc_hd__nand2_1 _07124_ (.A(_02101_),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__nand2_1 _07125_ (.A(_02003_),
    .B(_02082_),
    .Y(_02105_));
 sky130_fd_sc_hd__or3_1 _07126_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02079_),
    .C(_02099_),
    .X(_02106_));
 sky130_fd_sc_hd__nand2_1 _07127_ (.A(net3258),
    .B(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__o31a_1 _07128_ (.A1(_02099_),
    .A2(_02104_),
    .A3(_02105_),
    .B1(_02107_),
    .X(_02108_));
 sky130_fd_sc_hd__o21ai_1 _07129_ (.A1(_01997_),
    .A2(_02108_),
    .B1(_00614_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_1 _07130_ (.A(_01446_),
    .B(_02082_),
    .Y(_02109_));
 sky130_fd_sc_hd__nand2_1 _07131_ (.A(net3732),
    .B(_02106_),
    .Y(_02110_));
 sky130_fd_sc_hd__o31a_1 _07132_ (.A1(_02099_),
    .A2(_02104_),
    .A3(_02109_),
    .B1(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__o21ai_1 _07133_ (.A1(_01997_),
    .A2(_02111_),
    .B1(_01481_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__nand2_1 _07134_ (.A(_00551_),
    .B(_02082_),
    .Y(_02112_));
 sky130_fd_sc_hd__nand2_1 _07135_ (.A(net3593),
    .B(_02106_),
    .Y(_02113_));
 sky130_fd_sc_hd__o31a_1 _07136_ (.A1(_02099_),
    .A2(_02104_),
    .A3(_02112_),
    .B1(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__o21ai_1 _07137_ (.A1(_01997_),
    .A2(_02114_),
    .B1(_01912_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__nand2_1 _07138_ (.A(_01452_),
    .B(_02082_),
    .Y(_02115_));
 sky130_fd_sc_hd__nand2_1 _07139_ (.A(net3353),
    .B(_02106_),
    .Y(_02116_));
 sky130_fd_sc_hd__o31a_1 _07140_ (.A1(_02099_),
    .A2(_02104_),
    .A3(_02115_),
    .B1(_02116_),
    .X(_02117_));
 sky130_fd_sc_hd__buf_4 _07141_ (.A(_00226_),
    .X(_02118_));
 sky130_fd_sc_hd__o21ai_1 _07142_ (.A1(_01997_),
    .A2(_02117_),
    .B1(_02118_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _07143_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02079_),
    .Y(_02119_));
 sky130_fd_sc_hd__and3b_1 _07144_ (.A_N(_02089_),
    .B(_02088_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_02120_));
 sky130_fd_sc_hd__a21oi_4 _07145_ (.A1(_02119_),
    .A2(_02120_),
    .B1(_00267_),
    .Y(_02121_));
 sky130_fd_sc_hd__mux2_1 _07146_ (.A0(_02058_),
    .A1(net3427),
    .S(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__clkbuf_1 _07147_ (.A(_02122_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _07148_ (.A0(_02062_),
    .A1(net3450),
    .S(_02121_),
    .X(_02123_));
 sky130_fd_sc_hd__clkbuf_1 _07149_ (.A(_02123_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _07150_ (.A0(_02064_),
    .A1(net3553),
    .S(_02121_),
    .X(_02124_));
 sky130_fd_sc_hd__clkbuf_1 _07151_ (.A(_02124_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _07152_ (.A0(_01984_),
    .A1(net3615),
    .S(_02121_),
    .X(_02125_));
 sky130_fd_sc_hd__clkbuf_1 _07153_ (.A(_02125_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__clkbuf_4 _07154_ (.A(_00196_),
    .X(_02126_));
 sky130_fd_sc_hd__and4_1 _07155_ (.A(_02089_),
    .B(_02098_),
    .C(_02090_),
    .D(_02119_),
    .X(_02127_));
 sky130_fd_sc_hd__clkbuf_2 _07156_ (.A(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__nand2_1 _07157_ (.A(_02105_),
    .B(_02128_),
    .Y(_02129_));
 sky130_fd_sc_hd__or2_1 _07158_ (.A(net4097),
    .B(_02128_),
    .X(_02130_));
 sky130_fd_sc_hd__a31o_1 _07159_ (.A1(_02126_),
    .A2(_02129_),
    .A3(_02130_),
    .B1(_00603_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _07160_ (.A(_02109_),
    .B(_02128_),
    .Y(_02131_));
 sky130_fd_sc_hd__or2_1 _07161_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .B(_02128_),
    .X(_02132_));
 sky130_fd_sc_hd__clkbuf_8 _07162_ (.A(_00215_),
    .X(_02133_));
 sky130_fd_sc_hd__a31o_1 _07163_ (.A1(_02126_),
    .A2(_02131_),
    .A3(_02132_),
    .B1(_02133_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _07164_ (.A(_02112_),
    .B(_02128_),
    .Y(_02134_));
 sky130_fd_sc_hd__or2_1 _07165_ (.A(net4180),
    .B(_02128_),
    .X(_02135_));
 sky130_fd_sc_hd__a31o_1 _07166_ (.A1(_02126_),
    .A2(_02134_),
    .A3(_02135_),
    .B1(_00394_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _07167_ (.A(net4031),
    .B(_02128_),
    .Y(_02136_));
 sky130_fd_sc_hd__a211o_1 _07168_ (.A1(_02115_),
    .A2(_02128_),
    .B1(_02136_),
    .C1(_01471_),
    .X(_02137_));
 sky130_fd_sc_hd__nand2_1 _07169_ (.A(_02031_),
    .B(_02137_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _07170_ (.A1(_02089_),
    .A2(_02098_),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .A4(_02119_),
    .B1(_02034_),
    .X(_02138_));
 sky130_fd_sc_hd__mux2_1 _07171_ (.A0(net4073),
    .A1(_00692_),
    .S(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__clkbuf_1 _07172_ (.A(_02139_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _07173_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .A1(_00695_),
    .S(_02138_),
    .X(_02140_));
 sky130_fd_sc_hd__clkbuf_1 _07174_ (.A(_02140_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _07175_ (.A0(net3888),
    .A1(_00697_),
    .S(_02138_),
    .X(_02141_));
 sky130_fd_sc_hd__clkbuf_1 _07176_ (.A(_02141_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _07177_ (.A0(net3693),
    .A1(_02051_),
    .S(_02138_),
    .X(_02142_));
 sky130_fd_sc_hd__clkbuf_1 _07178_ (.A(_02142_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_1 _07179_ (.A(_02089_),
    .B(_02088_),
    .C(_02090_),
    .D(_02119_),
    .X(_02143_));
 sky130_fd_sc_hd__mux2_1 _07180_ (.A0(_01320_),
    .A1(_02105_),
    .S(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__clkbuf_8 _07181_ (.A(_00237_),
    .X(_02145_));
 sky130_fd_sc_hd__o21ai_1 _07182_ (.A1(_01997_),
    .A2(_02144_),
    .B1(_02145_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__clkbuf_4 _07183_ (.A(_00363_),
    .X(_02146_));
 sky130_fd_sc_hd__mux2_1 _07184_ (.A0(_01321_),
    .A1(_02109_),
    .S(_02143_),
    .X(_02147_));
 sky130_fd_sc_hd__o21ai_1 _07185_ (.A1(_02146_),
    .A2(_02147_),
    .B1(_01481_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__inv_2 _07186_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .Y(_02148_));
 sky130_fd_sc_hd__inv_2 _07187_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .Y(_02149_));
 sky130_fd_sc_hd__a31o_1 _07188_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .A2(_02149_),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_02150_));
 sky130_fd_sc_hd__or3b_1 _07189_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .B(_02150_),
    .C_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .X(_02151_));
 sky130_fd_sc_hd__o21ai_1 _07190_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ),
    .A2(_02148_),
    .B1(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__and2_1 _07191_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .B(_02150_),
    .X(_02153_));
 sky130_fd_sc_hd__mux4_1 _07192_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_02154_));
 sky130_fd_sc_hd__or2_1 _07193_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .B(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__mux2_1 _07194_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(_02156_));
 sky130_fd_sc_hd__inv_2 _07195_ (.A(net4030),
    .Y(_02157_));
 sky130_fd_sc_hd__mux2_1 _07196_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(_02158_));
 sky130_fd_sc_hd__inv_2 _07197_ (.A(net3848),
    .Y(_02159_));
 sky130_fd_sc_hd__a21o_1 _07198_ (.A1(_02157_),
    .A2(_02158_),
    .B1(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__a21o_1 _07199_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .A2(_02156_),
    .B1(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__mux4_1 _07200_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_02162_));
 sky130_fd_sc_hd__mux4_1 _07201_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(_02163_));
 sky130_fd_sc_hd__or2_1 _07202_ (.A(_02159_),
    .B(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__inv_2 _07203_ (.A(net3866),
    .Y(_02165_));
 sky130_fd_sc_hd__o211a_1 _07204_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .A2(_02162_),
    .B1(_02164_),
    .C1(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__a31oi_2 _07205_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ),
    .A2(_02155_),
    .A3(_02161_),
    .B1(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__and2b_1 _07206_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .X(_02168_));
 sky130_fd_sc_hd__a21bo_1 _07207_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_02169_));
 sky130_fd_sc_hd__mux2_1 _07208_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .X(_02170_));
 sky130_fd_sc_hd__o221a_1 _07209_ (.A1(_02168_),
    .A2(_02169_),
    .B1(_02170_),
    .B2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .X(_02171_));
 sky130_fd_sc_hd__inv_2 _07210_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .Y(_02172_));
 sky130_fd_sc_hd__mux4_1 _07211_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_02173_));
 sky130_fd_sc_hd__a21bo_1 _07212_ (.A1(_02172_),
    .A2(_02173_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(_02174_));
 sky130_fd_sc_hd__mux4_1 _07213_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_02175_));
 sky130_fd_sc_hd__mux4_1 _07214_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(_02176_));
 sky130_fd_sc_hd__mux2_1 _07215_ (.A0(_02175_),
    .A1(_02176_),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .X(_02177_));
 sky130_fd_sc_hd__o22a_4 _07216_ (.A1(_02171_),
    .A2(_02174_),
    .B1(_02177_),
    .B2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(_02178_));
 sky130_fd_sc_hd__mux2_1 _07217_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ),
    .S(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_1 _07218_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ),
    .S(_02178_),
    .X(_02180_));
 sky130_fd_sc_hd__inv_2 _07219_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .Y(_02181_));
 sky130_fd_sc_hd__mux4_1 _07220_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_02182_));
 sky130_fd_sc_hd__mux4_1 _07221_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_02183_));
 sky130_fd_sc_hd__mux2_1 _07222_ (.A0(_02182_),
    .A1(_02183_),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _07223_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(_02185_));
 sky130_fd_sc_hd__and2b_1 _07224_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .B(_02185_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _07225_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(_02187_));
 sky130_fd_sc_hd__a21bo_1 _07226_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .A2(_02187_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(_02188_));
 sky130_fd_sc_hd__mux4_1 _07227_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(_02189_));
 sky130_fd_sc_hd__o221a_1 _07228_ (.A1(_02186_),
    .A2(_02188_),
    .B1(_02189_),
    .B2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .X(_02190_));
 sky130_fd_sc_hd__a21o_2 _07229_ (.A1(_02181_),
    .A2(_02184_),
    .B1(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _07230_ (.A0(_02179_),
    .A1(_02180_),
    .S(_02191_),
    .X(_02192_));
 sky130_fd_sc_hd__and2_1 _07231_ (.A(_02167_),
    .B(_02192_),
    .X(_02193_));
 sky130_fd_sc_hd__a31o_1 _07232_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ),
    .A2(_02155_),
    .A3(_02161_),
    .B1(_02166_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _07233_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ),
    .S(_02178_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _07234_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ),
    .S(_02178_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _07235_ (.A0(_02195_),
    .A1(_02196_),
    .S(_02191_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _07236_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _07237_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_02199_));
 sky130_fd_sc_hd__or2b_1 _07238_ (.A(_02199_),
    .B_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(_02200_));
 sky130_fd_sc_hd__o211a_1 _07239_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_02198_),
    .B1(_02200_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _07240_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_02202_));
 sky130_fd_sc_hd__and2b_1 _07241_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .X(_02203_));
 sky130_fd_sc_hd__a21bo_1 _07242_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(_02204_));
 sky130_fd_sc_hd__inv_2 _07243_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .Y(_02205_));
 sky130_fd_sc_hd__o221a_1 _07244_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_02202_),
    .B1(_02203_),
    .B2(_02204_),
    .C1(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _07245_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_02207_));
 sky130_fd_sc_hd__or3b_1 _07246_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .C_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(_02208_));
 sky130_fd_sc_hd__o211a_1 _07247_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_02207_),
    .B1(_02208_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _07248_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_02210_));
 sky130_fd_sc_hd__inv_2 _07249_ (.A(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__mux2_1 _07250_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(_02212_));
 sky130_fd_sc_hd__nor2_1 _07251_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__a211o_1 _07252_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A2(_02211_),
    .B1(_02213_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(_02214_));
 sky130_fd_sc_hd__nand2_1 _07253_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .B(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__o32a_1 _07254_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .A2(_02201_),
    .A3(_02206_),
    .B1(_02209_),
    .B2(_02215_),
    .X(_02216_));
 sky130_fd_sc_hd__a21bo_1 _07255_ (.A1(_02194_),
    .A2(_02197_),
    .B1_N(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__mux2_1 _07256_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ),
    .S(_02178_),
    .X(_02218_));
 sky130_fd_sc_hd__mux2_1 _07257_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ),
    .S(_02178_),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _07258_ (.A0(_02218_),
    .A1(_02219_),
    .S(_02191_),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _07259_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ),
    .S(_02178_),
    .X(_02221_));
 sky130_fd_sc_hd__mux2_1 _07260_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ),
    .S(_02178_),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _07261_ (.A0(_02221_),
    .A1(_02222_),
    .S(_02191_),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _07262_ (.A0(_02220_),
    .A1(_02223_),
    .S(_02167_),
    .X(_02224_));
 sky130_fd_sc_hd__o221a_1 _07263_ (.A1(_02193_),
    .A2(_02217_),
    .B1(_02224_),
    .B2(_02216_),
    .C1(_01578_),
    .X(_02225_));
 sky130_fd_sc_hd__o2bb2a_4 _07264_ (.A1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .A2_N(_02152_),
    .B1(_02153_),
    .B2(_02225_),
    .X(_02226_));
 sky130_fd_sc_hd__buf_6 _07265_ (.A(_02226_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__mux2_1 _07266_ (.A0(_01324_),
    .A1(_02112_),
    .S(_02143_),
    .X(_02227_));
 sky130_fd_sc_hd__o21ai_1 _07267_ (.A1(_02146_),
    .A2(_02227_),
    .B1(_01912_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__buf_2 _07268_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .X(_02228_));
 sky130_fd_sc_hd__buf_2 _07269_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .X(_02229_));
 sky130_fd_sc_hd__mux4_1 _07270_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A2(_02228_),
    .A3(_02229_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .X(_02230_));
 sky130_fd_sc_hd__buf_2 _07271_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .X(_02231_));
 sky130_fd_sc_hd__clkbuf_4 _07272_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .X(_02232_));
 sky130_fd_sc_hd__clkbuf_4 _07273_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .X(_02233_));
 sky130_fd_sc_hd__clkbuf_4 _07274_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .X(_02234_));
 sky130_fd_sc_hd__mux4_1 _07275_ (.A0(_02231_),
    .A1(_02232_),
    .A2(_02233_),
    .A3(_02234_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _07276_ (.A0(_02230_),
    .A1(_02235_),
    .S(net3365),
    .X(_02236_));
 sky130_fd_sc_hd__clkbuf_1 _07277_ (.A(_02236_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ));
 sky130_fd_sc_hd__mux2_1 _07278_ (.A0(_01331_),
    .A1(_02115_),
    .S(_02143_),
    .X(_02237_));
 sky130_fd_sc_hd__o21ai_1 _07279_ (.A1(_02146_),
    .A2(_02237_),
    .B1(_02118_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a31o_1 _07280_ (.A1(_02149_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_02238_));
 sky130_fd_sc_hd__or3b_1 _07281_ (.A(_02238_),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .X(_02239_));
 sky130_fd_sc_hd__o21ai_1 _07282_ (.A1(_02148_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ),
    .B1(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__nand2_1 _07283_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .B(_02238_),
    .Y(_02241_));
 sky130_fd_sc_hd__mux2_1 _07284_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_02242_));
 sky130_fd_sc_hd__inv_2 _07285_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .Y(_02243_));
 sky130_fd_sc_hd__or3_1 _07286_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .C(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__o211ai_1 _07287_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_02242_),
    .B1(_02244_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .Y(_02245_));
 sky130_fd_sc_hd__mux2_1 _07288_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_1 _07289_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_02247_));
 sky130_fd_sc_hd__o21ba_1 _07290_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_02247_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_02248_));
 sky130_fd_sc_hd__o21ai_1 _07291_ (.A1(_02243_),
    .A2(_02246_),
    .B1(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hd__mux2_1 _07292_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_02250_));
 sky130_fd_sc_hd__or2_1 _07293_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .B(_02250_),
    .X(_02251_));
 sky130_fd_sc_hd__mux2_1 _07294_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_02252_));
 sky130_fd_sc_hd__o21a_1 _07295_ (.A1(_02243_),
    .A2(_02252_),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _07296_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _07297_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(_02255_));
 sky130_fd_sc_hd__o21ba_1 _07298_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A2(_02255_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(_02256_));
 sky130_fd_sc_hd__o21a_1 _07299_ (.A1(_02243_),
    .A2(_02254_),
    .B1(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__a211oi_1 _07300_ (.A1(_02251_),
    .A2(_02253_),
    .B1(_02257_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .Y(_02258_));
 sky130_fd_sc_hd__a31o_1 _07301_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .A2(_02245_),
    .A3(_02249_),
    .B1(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__inv_2 _07302_ (.A(net3690),
    .Y(_02260_));
 sky130_fd_sc_hd__mux4_1 _07303_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_02261_));
 sky130_fd_sc_hd__mux4_1 _07304_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_02262_));
 sky130_fd_sc_hd__inv_2 _07305_ (.A(net3687),
    .Y(_02263_));
 sky130_fd_sc_hd__mux2_1 _07306_ (.A0(_02261_),
    .A1(_02262_),
    .S(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__inv_2 _07307_ (.A(net4056),
    .Y(_02265_));
 sky130_fd_sc_hd__or2_1 _07308_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(_02266_));
 sky130_fd_sc_hd__o211a_1 _07309_ (.A1(_02265_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.half_q ),
    .B1(_02266_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_02267_));
 sky130_fd_sc_hd__inv_2 _07310_ (.A(net4092),
    .Y(_02268_));
 sky130_fd_sc_hd__mux2_1 _07311_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(_02269_));
 sky130_fd_sc_hd__a21o_1 _07312_ (.A1(_02268_),
    .A2(_02269_),
    .B1(_02263_),
    .X(_02270_));
 sky130_fd_sc_hd__mux4_1 _07313_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(_02271_));
 sky130_fd_sc_hd__or2_1 _07314_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .B(_02271_),
    .X(_02272_));
 sky130_fd_sc_hd__o211a_1 _07315_ (.A1(_02267_),
    .A2(_02270_),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ),
    .C1(_02272_),
    .X(_02273_));
 sky130_fd_sc_hd__a21oi_2 _07316_ (.A1(_02260_),
    .A2(_02264_),
    .B1(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__inv_2 _07317_ (.A(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hd__clkinv_2 _07318_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ),
    .Y(_02276_));
 sky130_fd_sc_hd__inv_2 _07319_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ),
    .Y(_02277_));
 sky130_fd_sc_hd__and2b_1 _07320_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .X(_02278_));
 sky130_fd_sc_hd__a21bo_1 _07321_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _07322_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .X(_02280_));
 sky130_fd_sc_hd__o221a_1 _07323_ (.A1(_02278_),
    .A2(_02279_),
    .B1(_02280_),
    .B2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .X(_02281_));
 sky130_fd_sc_hd__inv_2 _07324_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .Y(_02282_));
 sky130_fd_sc_hd__mux4_1 _07325_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_02283_));
 sky130_fd_sc_hd__a21bo_1 _07326_ (.A1(_02282_),
    .A2(_02283_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(_02284_));
 sky130_fd_sc_hd__mux4_1 _07327_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_02285_));
 sky130_fd_sc_hd__mux4_1 _07328_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _07329_ (.A0(_02285_),
    .A1(_02286_),
    .S(_02282_),
    .X(_02287_));
 sky130_fd_sc_hd__o22a_4 _07330_ (.A1(_02281_),
    .A2(_02284_),
    .B1(_02287_),
    .B2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _07331_ (.A0(_02276_),
    .A1(_02277_),
    .S(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__clkinv_2 _07332_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ),
    .Y(_02290_));
 sky130_fd_sc_hd__inv_2 _07333_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ),
    .Y(_02291_));
 sky130_fd_sc_hd__mux2_1 _07334_ (.A0(_02290_),
    .A1(_02291_),
    .S(_02288_),
    .X(_02292_));
 sky130_fd_sc_hd__inv_2 _07335_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .Y(_02293_));
 sky130_fd_sc_hd__mux4_1 _07336_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_02294_));
 sky130_fd_sc_hd__mux4_1 _07337_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _07338_ (.A0(_02294_),
    .A1(_02295_),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(_02296_));
 sky130_fd_sc_hd__mux4_1 _07339_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(_02297_));
 sky130_fd_sc_hd__mux2_1 _07340_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(_02298_));
 sky130_fd_sc_hd__and2b_1 _07341_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .B(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__mux2_1 _07342_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(_02300_));
 sky130_fd_sc_hd__a21bo_1 _07343_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .A2(_02300_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(_02301_));
 sky130_fd_sc_hd__o221a_1 _07344_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .A2(_02297_),
    .B1(_02299_),
    .B2(_02301_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .X(_02302_));
 sky130_fd_sc_hd__a21oi_2 _07345_ (.A1(_02293_),
    .A2(_02296_),
    .B1(_02302_),
    .Y(_02303_));
 sky130_fd_sc_hd__mux2_1 _07346_ (.A0(_02289_),
    .A1(_02292_),
    .S(_02303_),
    .X(_02304_));
 sky130_fd_sc_hd__inv_2 _07347_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ),
    .Y(_02305_));
 sky130_fd_sc_hd__nand2_1 _07348_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ),
    .B(_02288_),
    .Y(_02306_));
 sky130_fd_sc_hd__o211a_1 _07349_ (.A1(_02305_),
    .A2(_02288_),
    .B1(_02303_),
    .C1(_02306_),
    .X(_02307_));
 sky130_fd_sc_hd__mux2_1 _07350_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ),
    .S(_02288_),
    .X(_02308_));
 sky130_fd_sc_hd__o21bai_1 _07351_ (.A1(_02303_),
    .A2(_02308_),
    .B1_N(_02274_),
    .Y(_02309_));
 sky130_fd_sc_hd__o22a_1 _07352_ (.A1(_02275_),
    .A2(_02304_),
    .B1(_02307_),
    .B2(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _07353_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ),
    .S(_02288_),
    .X(_02311_));
 sky130_fd_sc_hd__mux2_1 _07354_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ),
    .S(_02288_),
    .X(_02312_));
 sky130_fd_sc_hd__mux2_1 _07355_ (.A0(_02311_),
    .A1(_02312_),
    .S(_02303_),
    .X(_02313_));
 sky130_fd_sc_hd__nand2_1 _07356_ (.A(_02274_),
    .B(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__mux2_1 _07357_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ),
    .S(_02288_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _07358_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ),
    .S(_02288_),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _07359_ (.A0(_02315_),
    .A1(_02316_),
    .S(_02303_),
    .X(_02317_));
 sky130_fd_sc_hd__a21oi_1 _07360_ (.A1(_02275_),
    .A2(_02317_),
    .B1(_02259_),
    .Y(_02318_));
 sky130_fd_sc_hd__a221o_2 _07361_ (.A1(_02259_),
    .A2(_02310_),
    .B1(_02314_),
    .B2(_02318_),
    .C1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ),
    .X(_02319_));
 sky130_fd_sc_hd__a22oi_4 _07362_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .A2(_02240_),
    .B1(_02241_),
    .B2(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hd__buf_6 _07363_ (.A(_02320_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__a41o_1 _07364_ (.A1(_02089_),
    .A2(_02088_),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .A4(_02119_),
    .B1(_02034_),
    .X(_02321_));
 sky130_fd_sc_hd__mux2_1 _07365_ (.A0(net4137),
    .A1(_00692_),
    .S(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__clkbuf_1 _07366_ (.A(_02322_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _07367_ (.A0(net4101),
    .A1(_00695_),
    .S(_02321_),
    .X(_02323_));
 sky130_fd_sc_hd__clkbuf_1 _07368_ (.A(_02323_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__buf_2 _07369_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ),
    .X(_02324_));
 sky130_fd_sc_hd__mux4_1 _07370_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(_02324_),
    .A2(_02231_),
    .A3(_02232_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(_02325_));
 sky130_fd_sc_hd__buf_2 _07371_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .X(_02326_));
 sky130_fd_sc_hd__mux4_1 _07372_ (.A0(_02326_),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(_02233_),
    .A3(_02234_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(_02327_));
 sky130_fd_sc_hd__mux2_1 _07373_ (.A0(_02325_),
    .A1(_02327_),
    .S(net3232),
    .X(_02328_));
 sky130_fd_sc_hd__clkbuf_1 _07374_ (.A(net3233),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ));
 sky130_fd_sc_hd__mux2_1 _07375_ (.A0(net3854),
    .A1(_00697_),
    .S(_02321_),
    .X(_02329_));
 sky130_fd_sc_hd__clkbuf_1 _07376_ (.A(_02329_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__a31o_1 _07377_ (.A1(_02149_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_02330_));
 sky130_fd_sc_hd__or3b_1 _07378_ (.A(_02330_),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .X(_02331_));
 sky130_fd_sc_hd__o21ai_1 _07379_ (.A1(_02148_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ),
    .B1(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__and2_1 _07380_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .B(_02330_),
    .X(_02333_));
 sky130_fd_sc_hd__mux2_1 _07381_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_02334_));
 sky130_fd_sc_hd__inv_2 _07382_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .Y(_02335_));
 sky130_fd_sc_hd__or3_1 _07383_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .C(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__o211ai_1 _07384_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_02334_),
    .B1(_02336_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .Y(_02337_));
 sky130_fd_sc_hd__mux2_1 _07385_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _07386_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_02339_));
 sky130_fd_sc_hd__o21ba_1 _07387_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_02339_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_02340_));
 sky130_fd_sc_hd__o21ai_1 _07388_ (.A1(_02335_),
    .A2(_02338_),
    .B1(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__mux2_1 _07389_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_02342_));
 sky130_fd_sc_hd__or2_1 _07390_ (.A(_02335_),
    .B(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__mux2_1 _07391_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_02344_));
 sky130_fd_sc_hd__o21a_1 _07392_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_02344_),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_02345_));
 sky130_fd_sc_hd__mux2_1 _07393_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_02346_));
 sky130_fd_sc_hd__mux2_1 _07394_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(_02347_));
 sky130_fd_sc_hd__o21ba_1 _07395_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A2(_02347_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(_02348_));
 sky130_fd_sc_hd__o21a_1 _07396_ (.A1(_02335_),
    .A2(_02346_),
    .B1(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__a211oi_1 _07397_ (.A1(_02343_),
    .A2(_02345_),
    .B1(_02349_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .Y(_02350_));
 sky130_fd_sc_hd__a31o_1 _07398_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .A2(_02337_),
    .A3(_02341_),
    .B1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__mux2_1 _07399_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .X(_02352_));
 sky130_fd_sc_hd__and2b_1 _07400_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .X(_02353_));
 sky130_fd_sc_hd__a21bo_1 _07401_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_02354_));
 sky130_fd_sc_hd__o221a_1 _07402_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .A2(_02352_),
    .B1(_02353_),
    .B2(_02354_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .X(_02355_));
 sky130_fd_sc_hd__inv_2 _07403_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .Y(_02356_));
 sky130_fd_sc_hd__mux4_1 _07404_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_02357_));
 sky130_fd_sc_hd__a21bo_1 _07405_ (.A1(_02356_),
    .A2(_02357_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .X(_02358_));
 sky130_fd_sc_hd__mux4_1 _07406_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_02359_));
 sky130_fd_sc_hd__mux4_1 _07407_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .X(_02360_));
 sky130_fd_sc_hd__mux2_1 _07408_ (.A0(_02359_),
    .A1(_02360_),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .X(_02361_));
 sky130_fd_sc_hd__o22a_4 _07409_ (.A1(_02355_),
    .A2(_02358_),
    .B1(_02361_),
    .B2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _07410_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ),
    .S(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__mux2_1 _07411_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ),
    .S(_02362_),
    .X(_02364_));
 sky130_fd_sc_hd__inv_2 _07412_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .Y(_02365_));
 sky130_fd_sc_hd__mux4_1 _07413_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_02366_));
 sky130_fd_sc_hd__mux4_1 _07414_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_02367_));
 sky130_fd_sc_hd__mux2_1 _07415_ (.A0(_02366_),
    .A1(_02367_),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_1 _07416_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(_02369_));
 sky130_fd_sc_hd__and2b_1 _07417_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .B(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__mux2_1 _07418_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(_02371_));
 sky130_fd_sc_hd__a21bo_1 _07419_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .A2(_02371_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(_02372_));
 sky130_fd_sc_hd__mux4_1 _07420_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(_02373_));
 sky130_fd_sc_hd__o221a_1 _07421_ (.A1(_02370_),
    .A2(_02372_),
    .B1(_02373_),
    .B2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .X(_02374_));
 sky130_fd_sc_hd__a21o_1 _07422_ (.A1(_02365_),
    .A2(_02368_),
    .B1(_02374_),
    .X(_02375_));
 sky130_fd_sc_hd__mux2_1 _07423_ (.A0(_02363_),
    .A1(_02364_),
    .S(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__mux2_1 _07424_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ),
    .S(_02362_),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _07425_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ),
    .S(_02362_),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _07426_ (.A0(_02377_),
    .A1(_02378_),
    .S(_02375_),
    .X(_02379_));
 sky130_fd_sc_hd__inv_2 _07427_ (.A(net3781),
    .Y(_02380_));
 sky130_fd_sc_hd__mux4_1 _07428_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_02381_));
 sky130_fd_sc_hd__mux4_1 _07429_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_02382_));
 sky130_fd_sc_hd__mux2_1 _07430_ (.A0(_02381_),
    .A1(_02382_),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .X(_02383_));
 sky130_fd_sc_hd__inv_2 _07431_ (.A(net4156),
    .Y(_02384_));
 sky130_fd_sc_hd__inv_2 _07432_ (.A(net3800),
    .Y(_02385_));
 sky130_fd_sc_hd__or2_1 _07433_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(_02386_));
 sky130_fd_sc_hd__o211a_1 _07434_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .A2(_02384_),
    .B1(_02385_),
    .C1(_02386_),
    .X(_02387_));
 sky130_fd_sc_hd__mux2_1 _07435_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(_02388_));
 sky130_fd_sc_hd__inv_2 _07436_ (.A(net3807),
    .Y(_02389_));
 sky130_fd_sc_hd__a21o_1 _07437_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .A2(_02388_),
    .B1(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__mux4_1 _07438_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(_02391_));
 sky130_fd_sc_hd__or2_1 _07439_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .B(_02391_),
    .X(_02392_));
 sky130_fd_sc_hd__o211a_1 _07440_ (.A1(_02387_),
    .A2(_02390_),
    .B1(_02392_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ),
    .X(_02393_));
 sky130_fd_sc_hd__a21oi_2 _07441_ (.A1(_02380_),
    .A2(_02383_),
    .B1(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__mux2_1 _07442_ (.A0(_02376_),
    .A1(_02379_),
    .S(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _07443_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ),
    .S(_02362_),
    .X(_02396_));
 sky130_fd_sc_hd__mux2_1 _07444_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ),
    .S(_02362_),
    .X(_02397_));
 sky130_fd_sc_hd__mux2_1 _07445_ (.A0(_02396_),
    .A1(_02397_),
    .S(_02375_),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _07446_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ),
    .S(_02362_),
    .X(_02399_));
 sky130_fd_sc_hd__or2_1 _07447_ (.A(_02375_),
    .B(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__clkinv_2 _07448_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ),
    .Y(_02401_));
 sky130_fd_sc_hd__clkinv_2 _07449_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ),
    .Y(_02402_));
 sky130_fd_sc_hd__mux2_1 _07450_ (.A0(_02401_),
    .A1(_02402_),
    .S(_02362_),
    .X(_02403_));
 sky130_fd_sc_hd__a21oi_1 _07451_ (.A1(_02375_),
    .A2(_02403_),
    .B1(_02394_),
    .Y(_02404_));
 sky130_fd_sc_hd__a31oi_2 _07452_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .A2(_02337_),
    .A3(_02341_),
    .B1(_02350_),
    .Y(_02405_));
 sky130_fd_sc_hd__a221o_1 _07453_ (.A1(_02394_),
    .A2(_02398_),
    .B1(_02400_),
    .B2(_02404_),
    .C1(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__o211a_2 _07454_ (.A1(_02351_),
    .A2(_02395_),
    .B1(_02406_),
    .C1(_01578_),
    .X(_02407_));
 sky130_fd_sc_hd__o2bb2a_4 _07455_ (.A1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .A2_N(_02332_),
    .B1(_02333_),
    .B2(_02407_),
    .X(_02408_));
 sky130_fd_sc_hd__buf_6 _07456_ (.A(_02408_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__mux2_1 _07457_ (.A0(net4011),
    .A1(_02051_),
    .S(_02321_),
    .X(_02409_));
 sky130_fd_sc_hd__clkbuf_1 _07458_ (.A(_02409_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__mux4_1 _07459_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A1(_02324_),
    .A2(_02326_),
    .A3(_02229_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .X(_02410_));
 sky130_fd_sc_hd__mux4_1 _07460_ (.A0(_02228_),
    .A1(_02232_),
    .A2(_02233_),
    .A3(_02234_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .X(_02411_));
 sky130_fd_sc_hd__mux2_1 _07461_ (.A0(_02410_),
    .A1(_02411_),
    .S(net3156),
    .X(_02412_));
 sky130_fd_sc_hd__clkbuf_1 _07462_ (.A(_02412_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ));
 sky130_fd_sc_hd__inv_2 _07463_ (.A(_02080_),
    .Y(_02413_));
 sky130_fd_sc_hd__a31o_2 _07464_ (.A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .A2(_02101_),
    .A3(_02413_),
    .B1(_00522_),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _07465_ (.A0(net3966),
    .A1(_00692_),
    .S(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__clkbuf_1 _07466_ (.A(_02415_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__a31o_1 _07467_ (.A1(_02149_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(_02416_));
 sky130_fd_sc_hd__or3b_1 _07468_ (.A(_02416_),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .C_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .X(_02417_));
 sky130_fd_sc_hd__o21ai_1 _07469_ (.A1(_02148_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ),
    .B1(_02417_),
    .Y(_02418_));
 sky130_fd_sc_hd__nand2_1 _07470_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .B(_02416_),
    .Y(_02419_));
 sky130_fd_sc_hd__inv_2 _07471_ (.A(net3521),
    .Y(_02420_));
 sky130_fd_sc_hd__mux4_1 _07472_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_02421_));
 sky130_fd_sc_hd__mux4_1 _07473_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _07474_ (.A0(_02421_),
    .A1(_02422_),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .X(_02423_));
 sky130_fd_sc_hd__mux4_1 _07475_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(_02424_));
 sky130_fd_sc_hd__inv_2 _07476_ (.A(net3937),
    .Y(_02425_));
 sky130_fd_sc_hd__inv_2 _07477_ (.A(net3982),
    .Y(_02426_));
 sky130_fd_sc_hd__or2_1 _07478_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(_02427_));
 sky130_fd_sc_hd__o211a_1 _07479_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .A2(_02425_),
    .B1(_02426_),
    .C1(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _07480_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.half_q ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(_02429_));
 sky130_fd_sc_hd__inv_2 _07481_ (.A(net3548),
    .Y(_02430_));
 sky130_fd_sc_hd__a21o_1 _07482_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .A2(_02429_),
    .B1(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__o221a_1 _07483_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .A2(_02424_),
    .B1(_02428_),
    .B2(_02431_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ),
    .X(_02432_));
 sky130_fd_sc_hd__a21o_1 _07484_ (.A1(_02420_),
    .A2(_02423_),
    .B1(_02432_),
    .X(_02433_));
 sky130_fd_sc_hd__and2b_1 _07485_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .X(_02434_));
 sky130_fd_sc_hd__a21bo_1 _07486_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _07487_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .X(_02436_));
 sky130_fd_sc_hd__o221a_1 _07488_ (.A1(_02434_),
    .A2(_02435_),
    .B1(_02436_),
    .B2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .X(_02437_));
 sky130_fd_sc_hd__inv_2 _07489_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .Y(_02438_));
 sky130_fd_sc_hd__mux4_1 _07490_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_02439_));
 sky130_fd_sc_hd__a21bo_1 _07491_ (.A1(_02438_),
    .A2(_02439_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .X(_02440_));
 sky130_fd_sc_hd__mux4_1 _07492_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_02441_));
 sky130_fd_sc_hd__mux4_1 _07493_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _07494_ (.A0(_02441_),
    .A1(_02442_),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .X(_02443_));
 sky130_fd_sc_hd__o22a_4 _07495_ (.A1(_02437_),
    .A2(_02440_),
    .B1(_02443_),
    .B2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _07496_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ),
    .S(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _07497_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ),
    .S(_02444_),
    .X(_02446_));
 sky130_fd_sc_hd__inv_2 _07498_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .Y(_02447_));
 sky130_fd_sc_hd__mux4_1 _07499_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_02448_));
 sky130_fd_sc_hd__mux4_1 _07500_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _07501_ (.A0(_02448_),
    .A1(_02449_),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(_02450_));
 sky130_fd_sc_hd__mux4_1 _07502_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _07503_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(_02452_));
 sky130_fd_sc_hd__and2b_1 _07504_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .B(_02452_),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _07505_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(_02454_));
 sky130_fd_sc_hd__a21bo_1 _07506_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .A2(_02454_),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(_02455_));
 sky130_fd_sc_hd__o221a_1 _07507_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .A2(_02451_),
    .B1(_02453_),
    .B2(_02455_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .X(_02456_));
 sky130_fd_sc_hd__a21oi_4 _07508_ (.A1(_02447_),
    .A2(_02450_),
    .B1(_02456_),
    .Y(_02457_));
 sky130_fd_sc_hd__mux2_1 _07509_ (.A0(_02445_),
    .A1(_02446_),
    .S(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__and2b_1 _07510_ (.A_N(_02433_),
    .B(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _07511_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ),
    .S(_02444_),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _07512_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ),
    .S(_02444_),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _07513_ (.A0(_02460_),
    .A1(_02461_),
    .S(_02457_),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _07514_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _07515_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_02464_));
 sky130_fd_sc_hd__or2b_1 _07516_ (.A(_02464_),
    .B_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .X(_02465_));
 sky130_fd_sc_hd__o211a_1 _07517_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_02463_),
    .B1(_02465_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _07518_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_02467_));
 sky130_fd_sc_hd__and2b_1 _07519_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .X(_02468_));
 sky130_fd_sc_hd__a21bo_1 _07520_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .B1_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .X(_02469_));
 sky130_fd_sc_hd__inv_2 _07521_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .Y(_02470_));
 sky130_fd_sc_hd__o221a_1 _07522_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_02467_),
    .B1(_02468_),
    .B2(_02469_),
    .C1(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _07523_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_02472_));
 sky130_fd_sc_hd__or3b_1 _07524_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .C_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .X(_02473_));
 sky130_fd_sc_hd__o211a_1 _07525_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_02472_),
    .B1(_02473_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _07526_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_02475_));
 sky130_fd_sc_hd__inv_2 _07527_ (.A(_02475_),
    .Y(_02476_));
 sky130_fd_sc_hd__mux2_1 _07528_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .S(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(_02477_));
 sky130_fd_sc_hd__nor2_1 _07529_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .B(_02477_),
    .Y(_02478_));
 sky130_fd_sc_hd__a211o_1 _07530_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A2(_02476_),
    .B1(_02478_),
    .C1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(_02479_));
 sky130_fd_sc_hd__nand2_1 _07531_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__o32a_1 _07532_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .A2(_02466_),
    .A3(_02471_),
    .B1(_02474_),
    .B2(_02480_),
    .X(_02481_));
 sky130_fd_sc_hd__a21bo_1 _07533_ (.A1(_02433_),
    .A2(_02462_),
    .B1_N(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _07534_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ),
    .S(_02444_),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _07535_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ),
    .S(_02444_),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _07536_ (.A0(_02483_),
    .A1(_02484_),
    .S(_02457_),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _07537_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ),
    .S(_02444_),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _07538_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ),
    .S(_02444_),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _07539_ (.A0(_02486_),
    .A1(_02487_),
    .S(_02457_),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _07540_ (.A0(_02485_),
    .A1(_02488_),
    .S(_02433_),
    .X(_02489_));
 sky130_fd_sc_hd__o221ai_4 _07541_ (.A1(_02459_),
    .A2(_02482_),
    .B1(_02489_),
    .B2(_02481_),
    .C1(_01578_),
    .Y(_02490_));
 sky130_fd_sc_hd__a22oi_4 _07542_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .A2(_02418_),
    .B1(_02419_),
    .B2(_02490_),
    .Y(_02491_));
 sky130_fd_sc_hd__buf_6 _07543_ (.A(_02491_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__mux2_1 _07544_ (.A0(net3602),
    .A1(_00695_),
    .S(_02414_),
    .X(_02492_));
 sky130_fd_sc_hd__clkbuf_1 _07545_ (.A(_02492_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _07546_ (.A0(net3868),
    .A1(_00697_),
    .S(_02414_),
    .X(_02493_));
 sky130_fd_sc_hd__clkbuf_1 _07547_ (.A(_02493_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux4_1 _07548_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A1(_02324_),
    .A2(_02326_),
    .A3(_02229_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .X(_02494_));
 sky130_fd_sc_hd__mux4_1 _07549_ (.A0(_02228_),
    .A1(_02231_),
    .A2(_02233_),
    .A3(_02234_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _07550_ (.A0(_02494_),
    .A1(_02495_),
    .S(net3585),
    .X(_02496_));
 sky130_fd_sc_hd__clkbuf_1 _07551_ (.A(_02496_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ));
 sky130_fd_sc_hd__mux2_1 _07552_ (.A0(net3958),
    .A1(_02051_),
    .S(_02414_),
    .X(_02497_));
 sky130_fd_sc_hd__clkbuf_1 _07553_ (.A(_02497_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _07554_ (.A(_02079_),
    .B(_02103_),
    .X(_02498_));
 sky130_fd_sc_hd__o41a_2 _07555_ (.A1(_02089_),
    .A2(_02088_),
    .A3(_02090_),
    .A4(_02498_),
    .B1(_01497_),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _07556_ (.A0(_02058_),
    .A1(net3833),
    .S(_02499_),
    .X(_02500_));
 sky130_fd_sc_hd__clkbuf_1 _07557_ (.A(_02500_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _07558_ (.A0(_02062_),
    .A1(net3484),
    .S(_02499_),
    .X(_02501_));
 sky130_fd_sc_hd__clkbuf_1 _07559_ (.A(_02501_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _07560_ (.A0(_02064_),
    .A1(net3976),
    .S(_02499_),
    .X(_02502_));
 sky130_fd_sc_hd__clkbuf_1 _07561_ (.A(_02502_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _07562_ (.A0(_01984_),
    .A1(net3518),
    .S(_02499_),
    .X(_02503_));
 sky130_fd_sc_hd__clkbuf_1 _07563_ (.A(_02503_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _07564_ (.A(_02099_),
    .B(_02498_),
    .Y(_02504_));
 sky130_fd_sc_hd__mux2_1 _07565_ (.A0(_01406_),
    .A1(_02105_),
    .S(_02504_),
    .X(_02505_));
 sky130_fd_sc_hd__o21ai_1 _07566_ (.A1(_02146_),
    .A2(_02505_),
    .B1(_02145_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__nand2_1 _07567_ (.A(_02109_),
    .B(_02504_),
    .Y(_02506_));
 sky130_fd_sc_hd__or2_1 _07568_ (.A(net4125),
    .B(_02504_),
    .X(_02507_));
 sky130_fd_sc_hd__a31o_1 _07569_ (.A1(_02126_),
    .A2(_02506_),
    .A3(_02507_),
    .B1(_02133_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__mux2_1 _07570_ (.A0(_01413_),
    .A1(_02112_),
    .S(_02504_),
    .X(_02508_));
 sky130_fd_sc_hd__o21ai_1 _07571_ (.A1(_02146_),
    .A2(_02508_),
    .B1(_01912_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__mux2_1 _07572_ (.A0(_01411_),
    .A1(_02115_),
    .S(_02504_),
    .X(_02509_));
 sky130_fd_sc_hd__o21ai_1 _07573_ (.A1(_02146_),
    .A2(_02509_),
    .B1(_02118_),
    .Y(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3_1 _07574_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02101_),
    .C(_02120_),
    .X(_02510_));
 sky130_fd_sc_hd__nor2_1 _07575_ (.A(_01971_),
    .B(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__a221o_1 _07576_ (.A1(_01762_),
    .A2(_02510_),
    .B1(_02511_),
    .B2(net3295),
    .C1(_01766_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _07577_ (.A1(_01771_),
    .A2(_02510_),
    .B1(_02511_),
    .B2(net3219),
    .C1(_01772_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _07578_ (.A1(_01850_),
    .A2(_02510_),
    .B1(_02511_),
    .B2(net3379),
    .C1(_01973_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__mux4_1 _07579_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A2(_02228_),
    .A3(_02229_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .X(_02512_));
 sky130_fd_sc_hd__mux4_1 _07580_ (.A0(_02231_),
    .A1(_02232_),
    .A2(_02233_),
    .A3(_02234_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _07581_ (.A0(_02512_),
    .A1(_02513_),
    .S(net3705),
    .X(_02514_));
 sky130_fd_sc_hd__clkbuf_1 _07582_ (.A(_02514_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ));
 sky130_fd_sc_hd__mux4_1 _07583_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(_02324_),
    .A2(_02231_),
    .A3(_02232_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ),
    .X(_02515_));
 sky130_fd_sc_hd__mux4_1 _07584_ (.A0(_02326_),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(_02233_),
    .A3(_02234_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _07585_ (.A0(_02515_),
    .A1(_02516_),
    .S(net3720),
    .X(_02517_));
 sky130_fd_sc_hd__clkbuf_1 _07586_ (.A(_02517_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ));
 sky130_fd_sc_hd__mux4_1 _07587_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A1(_02324_),
    .A2(_02326_),
    .A3(_02229_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ),
    .X(_02518_));
 sky130_fd_sc_hd__mux4_1 _07588_ (.A0(_02228_),
    .A1(_02232_),
    .A2(_02233_),
    .A3(_02234_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _07589_ (.A0(_02518_),
    .A1(_02519_),
    .S(net3541),
    .X(_02520_));
 sky130_fd_sc_hd__clkbuf_1 _07590_ (.A(_02520_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ));
 sky130_fd_sc_hd__mux4_1 _07591_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A1(_02324_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A3(_02229_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ),
    .X(_02521_));
 sky130_fd_sc_hd__mux4_1 _07592_ (.A0(_02228_),
    .A1(_02231_),
    .A2(_02233_),
    .A3(_02234_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _07593_ (.A0(_02521_),
    .A1(_02522_),
    .S(net3160),
    .X(_02523_));
 sky130_fd_sc_hd__clkbuf_1 _07594_ (.A(net3161),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ));
 sky130_fd_sc_hd__and2_4 _07595_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.m[0] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.m[1] ),
    .X(_02524_));
 sky130_fd_sc_hd__buf_6 _07596_ (.A(_02524_),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _07597_ (.A0(_01859_),
    .A1(_02077_),
    .S(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__clkbuf_1 _07598_ (.A(_02526_),
    .X(_00015_));
 sky130_fd_sc_hd__mux4_1 _07599_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A3(_02229_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .X(_02527_));
 sky130_fd_sc_hd__mux4_1 _07600_ (.A0(_02231_),
    .A1(_02232_),
    .A2(_02233_),
    .A3(_02234_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _07601_ (.A0(_02527_),
    .A1(_02528_),
    .S(net3291),
    .X(_02529_));
 sky130_fd_sc_hd__clkbuf_1 _07602_ (.A(net3292),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ));
 sky130_fd_sc_hd__mux4_1 _07603_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(_02324_),
    .A2(_02231_),
    .A3(_02232_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(_02530_));
 sky130_fd_sc_hd__mux4_1 _07604_ (.A0(_02326_),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _07605_ (.A0(_02530_),
    .A1(_02531_),
    .S(net3331),
    .X(_02532_));
 sky130_fd_sc_hd__clkbuf_1 _07606_ (.A(net3332),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ));
 sky130_fd_sc_hd__nand3b_2 _07607_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .B(_01878_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.cfgd ),
    .Y(_02533_));
 sky130_fd_sc_hd__or3_1 _07608_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_02534_));
 sky130_fd_sc_hd__or2_1 _07609_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__clkbuf_2 _07610_ (.A(_02535_),
    .X(_02536_));
 sky130_fd_sc_hd__o21a_2 _07611_ (.A1(_02533_),
    .A2(_02536_),
    .B1(_02092_),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _07612_ (.A0(_02058_),
    .A1(net3499),
    .S(_02537_),
    .X(_02538_));
 sky130_fd_sc_hd__clkbuf_1 _07613_ (.A(_02538_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _07614_ (.A0(_02062_),
    .A1(net3440),
    .S(_02537_),
    .X(_02539_));
 sky130_fd_sc_hd__clkbuf_1 _07615_ (.A(_02539_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__inv_2 _07616_ (.A(net3717),
    .Y(_02540_));
 sky130_fd_sc_hd__mux4_1 _07617_ (.A0(_02326_),
    .A1(_02229_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A3(_02324_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .S1(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__mux4_1 _07618_ (.A0(_02228_),
    .A1(_02232_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ),
    .X(_02542_));
 sky130_fd_sc_hd__mux2_1 _07619_ (.A0(_02541_),
    .A1(_02542_),
    .S(net3681),
    .X(_02543_));
 sky130_fd_sc_hd__clkbuf_1 _07620_ (.A(_02543_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ));
 sky130_fd_sc_hd__mux2_1 _07621_ (.A0(_02064_),
    .A1(net3152),
    .S(_02537_),
    .X(_02544_));
 sky130_fd_sc_hd__clkbuf_1 _07622_ (.A(_02544_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _07623_ (.A0(_01984_),
    .A1(net3147),
    .S(_02537_),
    .X(_02545_));
 sky130_fd_sc_hd__clkbuf_1 _07624_ (.A(_02545_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__inv_2 _07625_ (.A(net3206),
    .Y(_02546_));
 sky130_fd_sc_hd__mux4_1 _07626_ (.A0(_02326_),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A3(_02324_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .S1(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__mux4_1 _07627_ (.A0(_02228_),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .S1(net3206),
    .X(_02548_));
 sky130_fd_sc_hd__mux2_1 _07628_ (.A0(_02547_),
    .A1(_02548_),
    .S(net3223),
    .X(_02549_));
 sky130_fd_sc_hd__clkbuf_1 _07629_ (.A(_02549_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ));
 sky130_fd_sc_hd__buf_2 _07630_ (.A(net3899),
    .X(_02550_));
 sky130_fd_sc_hd__clkbuf_2 _07631_ (.A(net3803),
    .X(_02551_));
 sky130_fd_sc_hd__inv_2 _07632_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .Y(_02552_));
 sky130_fd_sc_hd__or4_1 _07633_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_02551_),
    .C(_02552_),
    .D(_02533_),
    .X(_02553_));
 sky130_fd_sc_hd__o21a_2 _07634_ (.A1(_02550_),
    .A2(_02553_),
    .B1(_02092_),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _07635_ (.A0(_02058_),
    .A1(net3513),
    .S(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__clkbuf_1 _07636_ (.A(_02555_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _07637_ (.A0(_02062_),
    .A1(net3145),
    .S(_02554_),
    .X(_02556_));
 sky130_fd_sc_hd__clkbuf_1 _07638_ (.A(_02556_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _07639_ (.A0(_02064_),
    .A1(net3544),
    .S(_02554_),
    .X(_02557_));
 sky130_fd_sc_hd__clkbuf_1 _07640_ (.A(_02557_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__buf_4 _07641_ (.A(_00191_),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _07642_ (.A0(_02558_),
    .A1(net3639),
    .S(_02554_),
    .X(_02559_));
 sky130_fd_sc_hd__clkbuf_1 _07643_ (.A(_02559_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _07644_ (.A(_02550_),
    .Y(_02560_));
 sky130_fd_sc_hd__or3_2 _07645_ (.A(_02551_),
    .B(_02560_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_02561_));
 sky130_fd_sc_hd__and3b_2 _07646_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .B(_00311_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.cfgd ),
    .X(_02562_));
 sky130_fd_sc_hd__nand2_1 _07647_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_02534_),
    .Y(_02563_));
 sky130_fd_sc_hd__and2_1 _07648_ (.A(_02536_),
    .B(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__nand2_1 _07649_ (.A(_02562_),
    .B(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__nand2_2 _07650_ (.A(_02003_),
    .B(_02536_),
    .Y(_02566_));
 sky130_fd_sc_hd__or3_1 _07651_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_02533_),
    .C(_02561_),
    .X(_02567_));
 sky130_fd_sc_hd__nand2_1 _07652_ (.A(net3793),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__o31a_1 _07653_ (.A1(_02561_),
    .A2(_02565_),
    .A3(_02566_),
    .B1(_02568_),
    .X(_02569_));
 sky130_fd_sc_hd__o21ai_1 _07654_ (.A1(_02146_),
    .A2(_02569_),
    .B1(_02145_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_1 _07655_ (.A(_01446_),
    .B(_02536_),
    .Y(_02570_));
 sky130_fd_sc_hd__nand2_1 _07656_ (.A(net3719),
    .B(_02567_),
    .Y(_02571_));
 sky130_fd_sc_hd__o31a_1 _07657_ (.A1(_02561_),
    .A2(_02565_),
    .A3(_02570_),
    .B1(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__o21ai_1 _07658_ (.A1(_02146_),
    .A2(_02572_),
    .B1(_01481_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__buf_8 _07659_ (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[2] ),
    .X(_02573_));
 sky130_fd_sc_hd__nand2_1 _07660_ (.A(_02573_),
    .B(_02536_),
    .Y(_02574_));
 sky130_fd_sc_hd__nand2_1 _07661_ (.A(net3768),
    .B(_02567_),
    .Y(_02575_));
 sky130_fd_sc_hd__o31a_1 _07662_ (.A1(_02561_),
    .A2(_02565_),
    .A3(_02574_),
    .B1(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__o21ai_1 _07663_ (.A1(_02146_),
    .A2(_02576_),
    .B1(_01912_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__nand2_2 _07664_ (.A(_01452_),
    .B(_02536_),
    .Y(_02577_));
 sky130_fd_sc_hd__nand2_1 _07665_ (.A(net3806),
    .B(_02567_),
    .Y(_02578_));
 sky130_fd_sc_hd__o31a_1 _07666_ (.A1(_02561_),
    .A2(_02565_),
    .A3(_02577_),
    .B1(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__o21ai_1 _07667_ (.A1(_02146_),
    .A2(_02579_),
    .B1(_02118_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _07668_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_02533_),
    .Y(_02580_));
 sky130_fd_sc_hd__and3b_2 _07669_ (.A_N(_02551_),
    .B(_02550_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_02581_));
 sky130_fd_sc_hd__a21oi_4 _07670_ (.A1(_02580_),
    .A2(_02581_),
    .B1(_00267_),
    .Y(_02582_));
 sky130_fd_sc_hd__mux2_1 _07671_ (.A0(_02058_),
    .A1(net3481),
    .S(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__clkbuf_1 _07672_ (.A(_02583_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _07673_ (.A0(_02062_),
    .A1(net3420),
    .S(_02582_),
    .X(_02584_));
 sky130_fd_sc_hd__clkbuf_1 _07674_ (.A(_02584_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _07675_ (.A0(_02064_),
    .A1(net3542),
    .S(_02582_),
    .X(_02585_));
 sky130_fd_sc_hd__clkbuf_1 _07676_ (.A(_02585_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _07677_ (.A0(_02558_),
    .A1(net3527),
    .S(_02582_),
    .X(_02586_));
 sky130_fd_sc_hd__clkbuf_1 _07678_ (.A(_02586_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4_1 _07679_ (.A(_02551_),
    .B(_02560_),
    .C(_02552_),
    .D(_02580_),
    .X(_02587_));
 sky130_fd_sc_hd__clkbuf_2 _07680_ (.A(_02587_),
    .X(_02588_));
 sky130_fd_sc_hd__nand2_1 _07681_ (.A(_02566_),
    .B(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__or2_1 _07682_ (.A(net4085),
    .B(_02588_),
    .X(_02590_));
 sky130_fd_sc_hd__a31o_1 _07683_ (.A1(_02126_),
    .A2(_02589_),
    .A3(_02590_),
    .B1(_00603_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _07684_ (.A(_02570_),
    .B(_02588_),
    .Y(_02591_));
 sky130_fd_sc_hd__or2_1 _07685_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .B(_02588_),
    .X(_02592_));
 sky130_fd_sc_hd__a31o_1 _07686_ (.A1(_02126_),
    .A2(_02591_),
    .A3(_02592_),
    .B1(_02133_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _07687_ (.A(_02574_),
    .B(_02588_),
    .Y(_02593_));
 sky130_fd_sc_hd__or2_1 _07688_ (.A(net4212),
    .B(_02588_),
    .X(_02594_));
 sky130_fd_sc_hd__a31o_1 _07689_ (.A1(_02126_),
    .A2(_02593_),
    .A3(_02594_),
    .B1(_00394_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _07690_ (.A(net4042),
    .B(_02588_),
    .Y(_02595_));
 sky130_fd_sc_hd__a211o_1 _07691_ (.A1(_02577_),
    .A2(_02588_),
    .B1(_02595_),
    .C1(_01471_),
    .X(_02596_));
 sky130_fd_sc_hd__nand2_1 _07692_ (.A(_02031_),
    .B(_02596_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__buf_4 _07693_ (.A(_00235_),
    .X(_02597_));
 sky130_fd_sc_hd__a41o_2 _07694_ (.A1(_02551_),
    .A2(_02560_),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .A4(_02580_),
    .B1(_02034_),
    .X(_02598_));
 sky130_fd_sc_hd__mux2_1 _07695_ (.A0(net4074),
    .A1(_02597_),
    .S(_02598_),
    .X(_02599_));
 sky130_fd_sc_hd__clkbuf_1 _07696_ (.A(_02599_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__buf_4 _07697_ (.A(_00292_),
    .X(_02600_));
 sky130_fd_sc_hd__mux2_1 _07698_ (.A0(net4201),
    .A1(_02600_),
    .S(_02598_),
    .X(_02601_));
 sky130_fd_sc_hd__clkbuf_1 _07699_ (.A(_02601_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__clkbuf_8 _07700_ (.A(_00188_),
    .X(_02602_));
 sky130_fd_sc_hd__mux2_1 _07701_ (.A0(net3986),
    .A1(_02602_),
    .S(_02598_),
    .X(_02603_));
 sky130_fd_sc_hd__clkbuf_1 _07702_ (.A(_02603_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _07703_ (.A0(net3874),
    .A1(_02051_),
    .S(_02598_),
    .X(_02604_));
 sky130_fd_sc_hd__clkbuf_1 _07704_ (.A(_02604_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__buf_2 _07705_ (.A(_01764_),
    .X(_02605_));
 sky130_fd_sc_hd__and4_1 _07706_ (.A(_02551_),
    .B(_02550_),
    .C(_02552_),
    .D(_02580_),
    .X(_02606_));
 sky130_fd_sc_hd__mux2_1 _07707_ (.A0(_01513_),
    .A1(_02566_),
    .S(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__o21ai_1 _07708_ (.A1(_02605_),
    .A2(_02607_),
    .B1(_02145_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _07709_ (.A0(_01516_),
    .A1(_02570_),
    .S(_02606_),
    .X(_02608_));
 sky130_fd_sc_hd__o21ai_1 _07710_ (.A1(_02605_),
    .A2(_02608_),
    .B1(_01481_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _07711_ (.A0(_01518_),
    .A1(_02574_),
    .S(_02606_),
    .X(_02609_));
 sky130_fd_sc_hd__o21ai_1 _07712_ (.A1(_02605_),
    .A2(_02609_),
    .B1(_01912_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _07713_ (.A0(_01508_),
    .A1(_02577_),
    .S(_02606_),
    .X(_02610_));
 sky130_fd_sc_hd__o21ai_1 _07714_ (.A1(_02605_),
    .A2(_02610_),
    .B1(_02118_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _07715_ (.A1(_02551_),
    .A2(_02550_),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .A4(_02580_),
    .B1(_02034_),
    .X(_02611_));
 sky130_fd_sc_hd__mux2_1 _07716_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .A1(_02597_),
    .S(_02611_),
    .X(_02612_));
 sky130_fd_sc_hd__clkbuf_1 _07717_ (.A(_02612_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _07718_ (.A0(net3955),
    .A1(_02600_),
    .S(_02611_),
    .X(_02613_));
 sky130_fd_sc_hd__clkbuf_1 _07719_ (.A(_02613_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _07720_ (.A0(net3782),
    .A1(_02602_),
    .S(_02611_),
    .X(_02614_));
 sky130_fd_sc_hd__clkbuf_1 _07721_ (.A(_02614_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _07722_ (.A0(net4128),
    .A1(_02051_),
    .S(_02611_),
    .X(_02615_));
 sky130_fd_sc_hd__clkbuf_1 _07723_ (.A(_02615_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _07724_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .Y(_02616_));
 sky130_fd_sc_hd__o31a_2 _07725_ (.A1(_02616_),
    .A2(_02533_),
    .A3(_02534_),
    .B1(_01489_),
    .X(_02617_));
 sky130_fd_sc_hd__mux2_1 _07726_ (.A0(_02058_),
    .A1(net3939),
    .S(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__clkbuf_1 _07727_ (.A(_02618_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _07728_ (.A0(_02062_),
    .A1(net3157),
    .S(_02617_),
    .X(_02619_));
 sky130_fd_sc_hd__clkbuf_1 _07729_ (.A(_02619_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _07730_ (.A0(_02064_),
    .A1(net3163),
    .S(_02617_),
    .X(_02620_));
 sky130_fd_sc_hd__clkbuf_1 _07731_ (.A(_02620_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _07732_ (.A0(_02558_),
    .A1(net3934),
    .S(_02617_),
    .X(_02621_));
 sky130_fd_sc_hd__clkbuf_1 _07733_ (.A(_02621_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _07734_ (.A(_02533_),
    .B(_02564_),
    .X(_02622_));
 sky130_fd_sc_hd__o41a_2 _07735_ (.A1(_02551_),
    .A2(_02550_),
    .A3(_02552_),
    .A4(_02622_),
    .B1(_01497_),
    .X(_02623_));
 sky130_fd_sc_hd__mux2_1 _07736_ (.A0(_02058_),
    .A1(net3909),
    .S(_02623_),
    .X(_02624_));
 sky130_fd_sc_hd__clkbuf_1 _07737_ (.A(_02624_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _07738_ (.A0(_02062_),
    .A1(net3555),
    .S(_02623_),
    .X(_02625_));
 sky130_fd_sc_hd__clkbuf_1 _07739_ (.A(_02625_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _07740_ (.A0(_02064_),
    .A1(net3865),
    .S(_02623_),
    .X(_02626_));
 sky130_fd_sc_hd__clkbuf_1 _07741_ (.A(_02626_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _07742_ (.A0(_02558_),
    .A1(net3459),
    .S(_02623_),
    .X(_02627_));
 sky130_fd_sc_hd__clkbuf_1 _07743_ (.A(_02627_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _07744_ (.A(_02561_),
    .B(_02622_),
    .Y(_02628_));
 sky130_fd_sc_hd__mux2_1 _07745_ (.A0(_01767_),
    .A1(_02566_),
    .S(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__o21ai_1 _07746_ (.A1(_02605_),
    .A2(_02629_),
    .B1(_02145_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__or2_1 _07747_ (.A(net4061),
    .B(_02628_),
    .X(_02630_));
 sky130_fd_sc_hd__nand2_1 _07748_ (.A(_02570_),
    .B(_02628_),
    .Y(_02631_));
 sky130_fd_sc_hd__a31o_1 _07749_ (.A1(_02126_),
    .A2(_02630_),
    .A3(_02631_),
    .B1(_02133_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__or2_1 _07750_ (.A(net3655),
    .B(_02628_),
    .X(_02632_));
 sky130_fd_sc_hd__nand2_1 _07751_ (.A(_02574_),
    .B(_02628_),
    .Y(_02633_));
 sky130_fd_sc_hd__buf_6 _07752_ (.A(_00221_),
    .X(_02634_));
 sky130_fd_sc_hd__a31o_1 _07753_ (.A1(_02126_),
    .A2(_02632_),
    .A3(_02633_),
    .B1(_02634_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__mux2_1 _07754_ (.A0(_01852_),
    .A1(_02577_),
    .S(_02628_),
    .X(_02635_));
 sky130_fd_sc_hd__o21ai_1 _07755_ (.A1(_02605_),
    .A2(_02635_),
    .B1(_02118_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3b_1 _07756_ (.A_N(_02564_),
    .B(_02581_),
    .C(_02562_),
    .X(_02636_));
 sky130_fd_sc_hd__buf_12 _07757_ (.A(_00249_),
    .X(_02637_));
 sky130_fd_sc_hd__a31oi_4 _07758_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .A2(_02562_),
    .A3(_02581_),
    .B1(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__a221o_1 _07759_ (.A1(_01762_),
    .A2(_02636_),
    .B1(_02638_),
    .B2(net3271),
    .C1(_01766_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _07760_ (.A1(_01771_),
    .A2(_02636_),
    .B1(_02638_),
    .B2(net3234),
    .C1(_01772_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _07761_ (.A1(_01850_),
    .A2(_02636_),
    .B1(_02638_),
    .B2(net3253),
    .C1(_01973_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__a22o_1 _07762_ (.A1(_01837_),
    .A2(_01841_),
    .B1(_01843_),
    .B2(_01845_),
    .X(_02639_));
 sky130_fd_sc_hd__and2_1 _07763_ (.A(_01858_),
    .B(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__and2_1 _07764_ (.A(_01858_),
    .B(_01577_),
    .X(_02641_));
 sky130_fd_sc_hd__mux2_1 _07765_ (.A0(_02640_),
    .A1(_02641_),
    .S(_01863_),
    .X(_02642_));
 sky130_fd_sc_hd__clkbuf_1 _07766_ (.A(_02642_),
    .X(_00008_));
 sky130_fd_sc_hd__clkbuf_4 _07767_ (.A(_00171_),
    .X(_02643_));
 sky130_fd_sc_hd__nand3b_2 _07768_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .C(_01415_),
    .Y(_02644_));
 sky130_fd_sc_hd__or3_1 _07769_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_02645_));
 sky130_fd_sc_hd__or2_1 _07770_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_02645_),
    .X(_02646_));
 sky130_fd_sc_hd__clkbuf_2 _07771_ (.A(_02646_),
    .X(_02647_));
 sky130_fd_sc_hd__o21a_2 _07772_ (.A1(_02644_),
    .A2(_02647_),
    .B1(_02092_),
    .X(_02648_));
 sky130_fd_sc_hd__mux2_1 _07773_ (.A0(_02643_),
    .A1(net3491),
    .S(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__clkbuf_1 _07774_ (.A(_02649_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__clkbuf_4 _07775_ (.A(_00184_),
    .X(_02650_));
 sky130_fd_sc_hd__mux2_1 _07776_ (.A0(_02650_),
    .A1(net3522),
    .S(_02648_),
    .X(_02651_));
 sky130_fd_sc_hd__clkbuf_1 _07777_ (.A(_02651_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__clkbuf_4 _07778_ (.A(_00551_),
    .X(_02652_));
 sky130_fd_sc_hd__mux2_1 _07779_ (.A0(_02652_),
    .A1(net3435),
    .S(_02648_),
    .X(_02653_));
 sky130_fd_sc_hd__clkbuf_1 _07780_ (.A(_02653_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _07781_ (.A0(_02558_),
    .A1(net3508),
    .S(_02648_),
    .X(_02654_));
 sky130_fd_sc_hd__clkbuf_1 _07782_ (.A(_02654_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _07783_ (.A(net4144),
    .X(_02655_));
 sky130_fd_sc_hd__clkbuf_2 _07784_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ),
    .X(_02656_));
 sky130_fd_sc_hd__inv_2 _07785_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .Y(_02657_));
 sky130_fd_sc_hd__or4_1 _07786_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_02656_),
    .C(_02657_),
    .D(_02644_),
    .X(_02658_));
 sky130_fd_sc_hd__o21a_2 _07787_ (.A1(_02655_),
    .A2(_02658_),
    .B1(_02092_),
    .X(_02659_));
 sky130_fd_sc_hd__mux2_1 _07788_ (.A0(_02643_),
    .A1(net3568),
    .S(_02659_),
    .X(_02660_));
 sky130_fd_sc_hd__clkbuf_1 _07789_ (.A(_02660_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _07790_ (.A0(_02650_),
    .A1(net3623),
    .S(_02659_),
    .X(_02661_));
 sky130_fd_sc_hd__clkbuf_1 _07791_ (.A(_02661_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _07792_ (.A0(_02652_),
    .A1(net3536),
    .S(_02659_),
    .X(_02662_));
 sky130_fd_sc_hd__clkbuf_1 _07793_ (.A(_02662_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _07794_ (.A0(_02558_),
    .A1(net3645),
    .S(_02659_),
    .X(_02663_));
 sky130_fd_sc_hd__clkbuf_1 _07795_ (.A(_02663_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _07796_ (.A(_02655_),
    .Y(_02664_));
 sky130_fd_sc_hd__or3_2 _07797_ (.A(_02656_),
    .B(_02664_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_02665_));
 sky130_fd_sc_hd__and3b_1 _07798_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .C(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ),
    .X(_02666_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07799_ (.A(_02666_),
    .X(_02667_));
 sky130_fd_sc_hd__nand2_1 _07800_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_02645_),
    .Y(_02668_));
 sky130_fd_sc_hd__and2_1 _07801_ (.A(_02647_),
    .B(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__nand2_1 _07802_ (.A(_02667_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__nand2_1 _07803_ (.A(_02003_),
    .B(_02647_),
    .Y(_02671_));
 sky130_fd_sc_hd__or3_1 _07804_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_02644_),
    .C(_02665_),
    .X(_02672_));
 sky130_fd_sc_hd__nand2_1 _07805_ (.A(net3772),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__o31a_1 _07806_ (.A1(_02665_),
    .A2(_02670_),
    .A3(_02671_),
    .B1(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__o21ai_1 _07807_ (.A1(_02605_),
    .A2(_02674_),
    .B1(_02145_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_1 _07808_ (.A(_00211_),
    .B(_02647_),
    .Y(_02675_));
 sky130_fd_sc_hd__nand2_1 _07809_ (.A(net3859),
    .B(_02672_),
    .Y(_02676_));
 sky130_fd_sc_hd__o31a_1 _07810_ (.A1(_02665_),
    .A2(_02670_),
    .A3(_02675_),
    .B1(_02676_),
    .X(_02677_));
 sky130_fd_sc_hd__o21ai_1 _07811_ (.A1(_02605_),
    .A2(_02677_),
    .B1(_01481_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__nand2_1 _07812_ (.A(_02573_),
    .B(_02647_),
    .Y(_02678_));
 sky130_fd_sc_hd__nand2_1 _07813_ (.A(net3731),
    .B(_02672_),
    .Y(_02679_));
 sky130_fd_sc_hd__o31a_1 _07814_ (.A1(_02665_),
    .A2(_02670_),
    .A3(_02678_),
    .B1(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__o21ai_1 _07815_ (.A1(_02605_),
    .A2(_02680_),
    .B1(_01912_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__nand2_2 _07816_ (.A(_00264_),
    .B(_02647_),
    .Y(_02681_));
 sky130_fd_sc_hd__nand2_1 _07817_ (.A(net3808),
    .B(_02672_),
    .Y(_02682_));
 sky130_fd_sc_hd__o31a_1 _07818_ (.A1(_02665_),
    .A2(_02670_),
    .A3(_02681_),
    .B1(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__o21ai_1 _07819_ (.A1(_02605_),
    .A2(_02683_),
    .B1(_02118_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _07820_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_02644_),
    .Y(_02684_));
 sky130_fd_sc_hd__and3b_1 _07821_ (.A_N(_02656_),
    .B(_02655_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_02685_));
 sky130_fd_sc_hd__buf_12 _07822_ (.A(_00180_),
    .X(_02686_));
 sky130_fd_sc_hd__a21oi_4 _07823_ (.A1(_02684_),
    .A2(_02685_),
    .B1(_02686_),
    .Y(_02687_));
 sky130_fd_sc_hd__mux2_1 _07824_ (.A0(_02643_),
    .A1(net3429),
    .S(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__clkbuf_1 _07825_ (.A(_02688_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _07826_ (.A0(_02650_),
    .A1(net3344),
    .S(_02687_),
    .X(_02689_));
 sky130_fd_sc_hd__clkbuf_1 _07827_ (.A(_02689_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _07828_ (.A0(_02652_),
    .A1(net3455),
    .S(_02687_),
    .X(_02690_));
 sky130_fd_sc_hd__clkbuf_1 _07829_ (.A(_02690_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _07830_ (.A0(_02558_),
    .A1(net3164),
    .S(_02687_),
    .X(_02691_));
 sky130_fd_sc_hd__clkbuf_1 _07831_ (.A(_02691_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4_1 _07832_ (.A(_02656_),
    .B(_02664_),
    .C(_02657_),
    .D(_02684_),
    .X(_02692_));
 sky130_fd_sc_hd__clkbuf_2 _07833_ (.A(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__nand2_1 _07834_ (.A(_02671_),
    .B(_02693_),
    .Y(_02694_));
 sky130_fd_sc_hd__or2_1 _07835_ (.A(net4126),
    .B(_02693_),
    .X(_02695_));
 sky130_fd_sc_hd__a31o_1 _07836_ (.A1(_02126_),
    .A2(_02694_),
    .A3(_02695_),
    .B1(_00603_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__clkbuf_4 _07837_ (.A(_00196_),
    .X(_02696_));
 sky130_fd_sc_hd__nand2_1 _07838_ (.A(_02675_),
    .B(_02693_),
    .Y(_02697_));
 sky130_fd_sc_hd__or2_1 _07839_ (.A(net4066),
    .B(_02693_),
    .X(_02698_));
 sky130_fd_sc_hd__a31o_1 _07840_ (.A1(_02696_),
    .A2(_02697_),
    .A3(_02698_),
    .B1(_02133_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _07841_ (.A(_02678_),
    .B(_02693_),
    .Y(_02699_));
 sky130_fd_sc_hd__or2_1 _07842_ (.A(net3992),
    .B(_02693_),
    .X(_02700_));
 sky130_fd_sc_hd__a31o_1 _07843_ (.A1(_02696_),
    .A2(_02699_),
    .A3(_02700_),
    .B1(_02634_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _07844_ (.A(net4034),
    .B(_02693_),
    .Y(_02701_));
 sky130_fd_sc_hd__a211o_1 _07845_ (.A1(_02681_),
    .A2(_02693_),
    .B1(_02701_),
    .C1(_01471_),
    .X(_02702_));
 sky130_fd_sc_hd__nand2_1 _07846_ (.A(_02031_),
    .B(_02702_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _07847_ (.A1(_02656_),
    .A2(_02664_),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .A4(_02684_),
    .B1(_02034_),
    .X(_02703_));
 sky130_fd_sc_hd__mux2_1 _07848_ (.A0(net4025),
    .A1(_02597_),
    .S(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__clkbuf_1 _07849_ (.A(_02704_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _07850_ (.A0(net4160),
    .A1(_02600_),
    .S(_02703_),
    .X(_02705_));
 sky130_fd_sc_hd__clkbuf_1 _07851_ (.A(_02705_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _07852_ (.A0(net3967),
    .A1(_02602_),
    .S(_02703_),
    .X(_02706_));
 sky130_fd_sc_hd__clkbuf_1 _07853_ (.A(_02706_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _07854_ (.A0(net3452),
    .A1(_02051_),
    .S(_02703_),
    .X(_02707_));
 sky130_fd_sc_hd__clkbuf_1 _07855_ (.A(_02707_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_1 _07856_ (.A(_02656_),
    .B(_02655_),
    .C(_02657_),
    .D(_02684_),
    .X(_02708_));
 sky130_fd_sc_hd__or2_1 _07857_ (.A(net4161),
    .B(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__nand2_1 _07858_ (.A(_02671_),
    .B(_02708_),
    .Y(_02710_));
 sky130_fd_sc_hd__buf_6 _07859_ (.A(_00208_),
    .X(_02711_));
 sky130_fd_sc_hd__a31o_1 _07860_ (.A1(_02696_),
    .A2(_02709_),
    .A3(_02710_),
    .B1(_02711_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__clkbuf_4 _07861_ (.A(_01764_),
    .X(_02712_));
 sky130_fd_sc_hd__mux2_1 _07862_ (.A0(_01621_),
    .A1(_02675_),
    .S(_02708_),
    .X(_02713_));
 sky130_fd_sc_hd__buf_6 _07863_ (.A(_00305_),
    .X(_02714_));
 sky130_fd_sc_hd__o21ai_1 _07864_ (.A1(_02712_),
    .A2(_02713_),
    .B1(_02714_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _07865_ (.A0(_01623_),
    .A1(_02678_),
    .S(_02708_),
    .X(_02715_));
 sky130_fd_sc_hd__o21ai_1 _07866_ (.A1(_02712_),
    .A2(_02715_),
    .B1(_01912_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _07867_ (.A0(_01629_),
    .A1(_02681_),
    .S(_02708_),
    .X(_02716_));
 sky130_fd_sc_hd__o21ai_1 _07868_ (.A1(_02712_),
    .A2(_02716_),
    .B1(_02118_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _07869_ (.A1(_02656_),
    .A2(_02655_),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .A4(_02684_),
    .B1(_02034_),
    .X(_02717_));
 sky130_fd_sc_hd__mux2_1 _07870_ (.A0(net4090),
    .A1(_02597_),
    .S(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__clkbuf_1 _07871_ (.A(_02718_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _07872_ (.A0(net4080),
    .A1(_02600_),
    .S(_02717_),
    .X(_02719_));
 sky130_fd_sc_hd__clkbuf_1 _07873_ (.A(_02719_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _07874_ (.A0(net3475),
    .A1(_02602_),
    .S(_02717_),
    .X(_02720_));
 sky130_fd_sc_hd__clkbuf_1 _07875_ (.A(_02720_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _07876_ (.A0(net3898),
    .A1(_02051_),
    .S(_02717_),
    .X(_02721_));
 sky130_fd_sc_hd__clkbuf_1 _07877_ (.A(_02721_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _07878_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .Y(_02722_));
 sky130_fd_sc_hd__o31a_2 _07879_ (.A1(_02722_),
    .A2(_02644_),
    .A3(_02645_),
    .B1(_01489_),
    .X(_02723_));
 sky130_fd_sc_hd__mux2_1 _07880_ (.A0(_02643_),
    .A1(net3722),
    .S(_02723_),
    .X(_02724_));
 sky130_fd_sc_hd__clkbuf_1 _07881_ (.A(_02724_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _07882_ (.A0(_02650_),
    .A1(net3676),
    .S(_02723_),
    .X(_02725_));
 sky130_fd_sc_hd__clkbuf_1 _07883_ (.A(_02725_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _07884_ (.A0(_02652_),
    .A1(net3852),
    .S(_02723_),
    .X(_02726_));
 sky130_fd_sc_hd__clkbuf_1 _07885_ (.A(_02726_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _07886_ (.A0(_02558_),
    .A1(net3949),
    .S(_02723_),
    .X(_02727_));
 sky130_fd_sc_hd__clkbuf_1 _07887_ (.A(_02727_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _07888_ (.A(_02644_),
    .B(_02669_),
    .X(_02728_));
 sky130_fd_sc_hd__o41a_2 _07889_ (.A1(_02656_),
    .A2(_02655_),
    .A3(_02657_),
    .A4(_02728_),
    .B1(_01497_),
    .X(_02729_));
 sky130_fd_sc_hd__mux2_1 _07890_ (.A0(_02643_),
    .A1(net3801),
    .S(_02729_),
    .X(_02730_));
 sky130_fd_sc_hd__clkbuf_1 _07891_ (.A(_02730_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _07892_ (.A0(_02650_),
    .A1(net3262),
    .S(_02729_),
    .X(_02731_));
 sky130_fd_sc_hd__clkbuf_1 _07893_ (.A(_02731_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _07894_ (.A0(_02652_),
    .A1(net3931),
    .S(_02729_),
    .X(_02732_));
 sky130_fd_sc_hd__clkbuf_1 _07895_ (.A(_02732_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _07896_ (.A0(_02558_),
    .A1(net3654),
    .S(_02729_),
    .X(_02733_));
 sky130_fd_sc_hd__clkbuf_1 _07897_ (.A(_02733_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _07898_ (.A(_02665_),
    .B(_02728_),
    .Y(_02734_));
 sky130_fd_sc_hd__nand2_1 _07899_ (.A(_02671_),
    .B(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__or2_1 _07900_ (.A(net3851),
    .B(_02734_),
    .X(_02736_));
 sky130_fd_sc_hd__a31o_1 _07901_ (.A1(_02696_),
    .A2(_02735_),
    .A3(_02736_),
    .B1(_02711_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__or2_1 _07902_ (.A(net4077),
    .B(_02734_),
    .X(_02737_));
 sky130_fd_sc_hd__nand2_1 _07903_ (.A(_02675_),
    .B(_02734_),
    .Y(_02738_));
 sky130_fd_sc_hd__a31o_1 _07904_ (.A1(_02696_),
    .A2(_02737_),
    .A3(_02738_),
    .B1(_02133_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__mux2_1 _07905_ (.A0(_01876_),
    .A1(_02678_),
    .S(_02734_),
    .X(_02739_));
 sky130_fd_sc_hd__buf_6 _07906_ (.A(_00250_),
    .X(_02740_));
 sky130_fd_sc_hd__o21ai_1 _07907_ (.A1(_02712_),
    .A2(_02739_),
    .B1(_02740_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__nor2_1 _07908_ (.A(net3798),
    .B(_02734_),
    .Y(_02741_));
 sky130_fd_sc_hd__a211o_1 _07909_ (.A1(_02681_),
    .A2(_02734_),
    .B1(_02741_),
    .C1(_01471_),
    .X(_02742_));
 sky130_fd_sc_hd__nand2_1 _07910_ (.A(_02031_),
    .B(_02742_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3_2 _07911_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_02667_),
    .C(_02685_),
    .X(_02743_));
 sky130_fd_sc_hd__nor2_1 _07912_ (.A(_01971_),
    .B(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__a221o_1 _07913_ (.A1(_01762_),
    .A2(_02743_),
    .B1(_02744_),
    .B2(net3155),
    .C1(_01766_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _07914_ (.A1(_01771_),
    .A2(_02743_),
    .B1(_02744_),
    .B2(net3231),
    .C1(_01772_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _07915_ (.A1(_01850_),
    .A2(_02743_),
    .B1(_02744_),
    .B2(net3181),
    .C1(_01973_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__mux4_1 _07916_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A3(_01585_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .X(_02745_));
 sky130_fd_sc_hd__mux4_1 _07917_ (.A0(_01587_),
    .A1(_01588_),
    .A2(_01589_),
    .A3(_01590_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .X(_02746_));
 sky130_fd_sc_hd__mux2_1 _07918_ (.A0(_02745_),
    .A1(_02746_),
    .S(net3197),
    .X(_02747_));
 sky130_fd_sc_hd__clkbuf_1 _07919_ (.A(net3198),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ));
 sky130_fd_sc_hd__mux4_1 _07920_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(_01676_),
    .A2(_01587_),
    .A3(_01588_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .S1(net3318),
    .X(_02748_));
 sky130_fd_sc_hd__mux4_1 _07921_ (.A0(_01678_),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .S1(net3318),
    .X(_02749_));
 sky130_fd_sc_hd__mux2_1 _07922_ (.A0(_02748_),
    .A1(_02749_),
    .S(net3466),
    .X(_02750_));
 sky130_fd_sc_hd__clkbuf_1 _07923_ (.A(_02750_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ));
 sky130_fd_sc_hd__inv_2 _07924_ (.A(net3668),
    .Y(_02751_));
 sky130_fd_sc_hd__mux4_1 _07925_ (.A0(_01678_),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A3(_01676_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .S1(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__mux4_1 _07926_ (.A0(_01584_),
    .A1(_01588_),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ),
    .X(_02753_));
 sky130_fd_sc_hd__mux2_1 _07927_ (.A0(_02752_),
    .A1(_02753_),
    .S(net3361),
    .X(_02754_));
 sky130_fd_sc_hd__clkbuf_1 _07928_ (.A(net3362),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ));
 sky130_fd_sc_hd__inv_2 _07929_ (.A(net3929),
    .Y(_02755_));
 sky130_fd_sc_hd__mux4_1 _07930_ (.A0(_01678_),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A3(_01676_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .S1(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__mux4_1 _07931_ (.A0(_01584_),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ),
    .X(_02757_));
 sky130_fd_sc_hd__mux2_1 _07932_ (.A0(_02756_),
    .A1(_02757_),
    .S(net3394),
    .X(_02758_));
 sky130_fd_sc_hd__clkbuf_1 _07933_ (.A(_02758_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ));
 sky130_fd_sc_hd__buf_6 _07934_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ),
    .X(_02759_));
 sky130_fd_sc_hd__a21oi_1 _07935_ (.A1(_01657_),
    .A2(_01662_),
    .B1(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__mux2_1 _07936_ (.A0(_02641_),
    .A1(_02760_),
    .S(_01863_),
    .X(_02761_));
 sky130_fd_sc_hd__clkbuf_1 _07937_ (.A(_02761_),
    .X(_00009_));
 sky130_fd_sc_hd__nand3b_2 _07938_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .C(_01878_),
    .Y(_02762_));
 sky130_fd_sc_hd__or3_1 _07939_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_02763_));
 sky130_fd_sc_hd__or2_1 _07940_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07941_ (.A(_02764_),
    .X(_02765_));
 sky130_fd_sc_hd__o21a_2 _07942_ (.A1(_02762_),
    .A2(_02765_),
    .B1(_02092_),
    .X(_02766_));
 sky130_fd_sc_hd__mux2_1 _07943_ (.A0(_02643_),
    .A1(net3439),
    .S(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__clkbuf_1 _07944_ (.A(_02767_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _07945_ (.A0(_02650_),
    .A1(net3500),
    .S(_02766_),
    .X(_02768_));
 sky130_fd_sc_hd__clkbuf_1 _07946_ (.A(_02768_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _07947_ (.A0(_02652_),
    .A1(net3458),
    .S(_02766_),
    .X(_02769_));
 sky130_fd_sc_hd__clkbuf_1 _07948_ (.A(_02769_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _07949_ (.A0(_02558_),
    .A1(net3359),
    .S(_02766_),
    .X(_02770_));
 sky130_fd_sc_hd__clkbuf_1 _07950_ (.A(_02770_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _07951_ (.A(net4146),
    .X(_02771_));
 sky130_fd_sc_hd__clkbuf_2 _07952_ (.A(net4198),
    .X(_02772_));
 sky130_fd_sc_hd__inv_2 _07953_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .Y(_02773_));
 sky130_fd_sc_hd__or4_1 _07954_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_02772_),
    .C(_02773_),
    .D(_02762_),
    .X(_02774_));
 sky130_fd_sc_hd__o21a_2 _07955_ (.A1(_02771_),
    .A2(_02774_),
    .B1(_02092_),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_1 _07956_ (.A0(_02643_),
    .A1(net3296),
    .S(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__clkbuf_1 _07957_ (.A(_02776_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _07958_ (.A0(_02650_),
    .A1(net3501),
    .S(_02775_),
    .X(_02777_));
 sky130_fd_sc_hd__clkbuf_1 _07959_ (.A(_02777_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _07960_ (.A0(_02652_),
    .A1(net3579),
    .S(_02775_),
    .X(_02778_));
 sky130_fd_sc_hd__clkbuf_1 _07961_ (.A(_02778_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__clkbuf_4 _07962_ (.A(_00191_),
    .X(_02779_));
 sky130_fd_sc_hd__mux2_1 _07963_ (.A0(_02779_),
    .A1(net3461),
    .S(_02775_),
    .X(_02780_));
 sky130_fd_sc_hd__clkbuf_1 _07964_ (.A(_02780_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _07965_ (.A(_02771_),
    .Y(_02781_));
 sky130_fd_sc_hd__or3_2 _07966_ (.A(_02772_),
    .B(_02781_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_02782_));
 sky130_fd_sc_hd__and3b_1 _07967_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .C(_01415_),
    .X(_02783_));
 sky130_fd_sc_hd__nand2_1 _07968_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_02763_),
    .Y(_02784_));
 sky130_fd_sc_hd__and2_1 _07969_ (.A(_02765_),
    .B(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__nand2_1 _07970_ (.A(_02783_),
    .B(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__nand2_1 _07971_ (.A(_02003_),
    .B(_02765_),
    .Y(_02787_));
 sky130_fd_sc_hd__or3_1 _07972_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_02762_),
    .C(_02782_),
    .X(_02788_));
 sky130_fd_sc_hd__nand2_1 _07973_ (.A(net3627),
    .B(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__o31a_1 _07974_ (.A1(_02782_),
    .A2(_02786_),
    .A3(_02787_),
    .B1(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__o21ai_1 _07975_ (.A1(_02712_),
    .A2(_02790_),
    .B1(_02145_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_1 _07976_ (.A(_00211_),
    .B(_02765_),
    .Y(_02791_));
 sky130_fd_sc_hd__nand2_1 _07977_ (.A(net3590),
    .B(_02788_),
    .Y(_02792_));
 sky130_fd_sc_hd__o31a_1 _07978_ (.A1(_02782_),
    .A2(_02786_),
    .A3(_02791_),
    .B1(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__o21ai_1 _07979_ (.A1(_02712_),
    .A2(_02793_),
    .B1(_02714_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__nand2_1 _07980_ (.A(_02573_),
    .B(_02765_),
    .Y(_02794_));
 sky130_fd_sc_hd__nand2_1 _07981_ (.A(net3571),
    .B(_02788_),
    .Y(_02795_));
 sky130_fd_sc_hd__o31a_1 _07982_ (.A1(_02782_),
    .A2(_02786_),
    .A3(_02794_),
    .B1(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__o21ai_1 _07983_ (.A1(_02712_),
    .A2(_02796_),
    .B1(_02740_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__nand2_1 _07984_ (.A(_00264_),
    .B(_02765_),
    .Y(_02797_));
 sky130_fd_sc_hd__nand2_1 _07985_ (.A(net3736),
    .B(_02788_),
    .Y(_02798_));
 sky130_fd_sc_hd__o31a_1 _07986_ (.A1(_02782_),
    .A2(_02786_),
    .A3(_02797_),
    .B1(_02798_),
    .X(_02799_));
 sky130_fd_sc_hd__o21ai_1 _07987_ (.A1(_02712_),
    .A2(_02799_),
    .B1(_02118_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _07988_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_02762_),
    .Y(_02800_));
 sky130_fd_sc_hd__and3b_1 _07989_ (.A_N(_02772_),
    .B(_02771_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_02801_));
 sky130_fd_sc_hd__a21oi_4 _07990_ (.A1(_02800_),
    .A2(_02801_),
    .B1(_02686_),
    .Y(_02802_));
 sky130_fd_sc_hd__mux2_1 _07991_ (.A0(_02643_),
    .A1(net3437),
    .S(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__clkbuf_1 _07992_ (.A(_02803_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _07993_ (.A0(_02650_),
    .A1(net3324),
    .S(_02802_),
    .X(_02804_));
 sky130_fd_sc_hd__clkbuf_1 _07994_ (.A(_02804_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _07995_ (.A0(_02652_),
    .A1(net3345),
    .S(_02802_),
    .X(_02805_));
 sky130_fd_sc_hd__clkbuf_1 _07996_ (.A(_02805_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _07997_ (.A0(_02779_),
    .A1(net3326),
    .S(_02802_),
    .X(_02806_));
 sky130_fd_sc_hd__clkbuf_1 _07998_ (.A(_02806_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__mux4_1 _07999_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A3(_02229_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .X(_02807_));
 sky130_fd_sc_hd__mux4_1 _08000_ (.A0(_02231_),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _08001_ (.A0(_02807_),
    .A1(_02808_),
    .S(net3442),
    .X(_02809_));
 sky130_fd_sc_hd__clkbuf_1 _08002_ (.A(_02809_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ));
 sky130_fd_sc_hd__and4_1 _08003_ (.A(_02772_),
    .B(_02781_),
    .C(_02773_),
    .D(_02800_),
    .X(_02810_));
 sky130_fd_sc_hd__clkbuf_2 _08004_ (.A(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__nand2_1 _08005_ (.A(_02787_),
    .B(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__or2_1 _08006_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .B(_02811_),
    .X(_02813_));
 sky130_fd_sc_hd__a31o_1 _08007_ (.A1(_02696_),
    .A2(_02812_),
    .A3(_02813_),
    .B1(_02711_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _08008_ (.A(_02791_),
    .B(_02811_),
    .Y(_02814_));
 sky130_fd_sc_hd__or2_1 _08009_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .B(_02811_),
    .X(_02815_));
 sky130_fd_sc_hd__a31o_1 _08010_ (.A1(_02696_),
    .A2(_02814_),
    .A3(_02815_),
    .B1(_02133_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _08011_ (.A(_02794_),
    .B(_02811_),
    .Y(_02816_));
 sky130_fd_sc_hd__or2_1 _08012_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .B(_02811_),
    .X(_02817_));
 sky130_fd_sc_hd__a31o_1 _08013_ (.A1(_02696_),
    .A2(_02816_),
    .A3(_02817_),
    .B1(_02634_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__mux4_1 _08014_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ),
    .A2(_02231_),
    .A3(_02232_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .S1(net3617),
    .X(_02818_));
 sky130_fd_sc_hd__mux4_1 _08015_ (.A0(_02326_),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .S1(net3617),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_1 _08016_ (.A0(_02818_),
    .A1(_02819_),
    .S(net3380),
    .X(_02820_));
 sky130_fd_sc_hd__clkbuf_1 _08017_ (.A(_02820_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ));
 sky130_fd_sc_hd__nor2_1 _08018_ (.A(net4082),
    .B(_02811_),
    .Y(_02821_));
 sky130_fd_sc_hd__a211o_1 _08019_ (.A1(_02797_),
    .A2(_02811_),
    .B1(_02821_),
    .C1(_01471_),
    .X(_02822_));
 sky130_fd_sc_hd__nand2_1 _08020_ (.A(_02031_),
    .B(_02822_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _08021_ (.A1(_02772_),
    .A2(_02781_),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .A4(_02800_),
    .B1(_02034_),
    .X(_02823_));
 sky130_fd_sc_hd__mux2_1 _08022_ (.A0(net4050),
    .A1(_02597_),
    .S(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__clkbuf_1 _08023_ (.A(_02824_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux4_1 _08024_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A3(_02229_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .X(_02825_));
 sky130_fd_sc_hd__mux4_1 _08025_ (.A0(_02228_),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _08026_ (.A0(_02825_),
    .A1(_02826_),
    .S(net3605),
    .X(_02827_));
 sky130_fd_sc_hd__clkbuf_1 _08027_ (.A(_02827_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ));
 sky130_fd_sc_hd__mux2_1 _08028_ (.A0(net4204),
    .A1(_02600_),
    .S(_02823_),
    .X(_02828_));
 sky130_fd_sc_hd__clkbuf_1 _08029_ (.A(_02828_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _08030_ (.A0(net3860),
    .A1(_02602_),
    .S(_02823_),
    .X(_02829_));
 sky130_fd_sc_hd__clkbuf_1 _08031_ (.A(_02829_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__inv_2 _08032_ (.A(net3387),
    .Y(_02830_));
 sky130_fd_sc_hd__mux4_1 _08033_ (.A0(_02326_),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A3(_02324_),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .S1(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__mux4_1 _08034_ (.A0(_02228_),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .S1(net3387),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _08035_ (.A0(_02831_),
    .A1(_02832_),
    .S(net3523),
    .X(_02833_));
 sky130_fd_sc_hd__clkbuf_1 _08036_ (.A(_02833_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ));
 sky130_fd_sc_hd__mux2_1 _08037_ (.A0(net3876),
    .A1(_02051_),
    .S(_02823_),
    .X(_02834_));
 sky130_fd_sc_hd__clkbuf_1 _08038_ (.A(_02834_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_1 _08039_ (.A(_02772_),
    .B(_02771_),
    .C(_02773_),
    .D(_02800_),
    .X(_02835_));
 sky130_fd_sc_hd__mux2_1 _08040_ (.A0(_01691_),
    .A1(_02787_),
    .S(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__o21ai_1 _08041_ (.A1(_02712_),
    .A2(_02836_),
    .B1(_02145_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _08042_ (.A0(_01692_),
    .A1(_02791_),
    .S(_02835_),
    .X(_02837_));
 sky130_fd_sc_hd__o21ai_1 _08043_ (.A1(_02712_),
    .A2(_02837_),
    .B1(_02714_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__clkbuf_4 _08044_ (.A(_01764_),
    .X(_02838_));
 sky130_fd_sc_hd__mux2_1 _08045_ (.A0(_01696_),
    .A1(_02794_),
    .S(_02835_),
    .X(_02839_));
 sky130_fd_sc_hd__o21ai_1 _08046_ (.A1(_02838_),
    .A2(_02839_),
    .B1(_02740_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _08047_ (.A0(_01686_),
    .A1(_02797_),
    .S(_02835_),
    .X(_02840_));
 sky130_fd_sc_hd__o21ai_1 _08048_ (.A1(_02838_),
    .A2(_02840_),
    .B1(_02118_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _08049_ (.A1(_02772_),
    .A2(_02771_),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .A4(_02800_),
    .B1(_02034_),
    .X(_02841_));
 sky130_fd_sc_hd__mux2_1 _08050_ (.A0(net4177),
    .A1(_02597_),
    .S(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_1 _08051_ (.A(_02842_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _08052_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .A1(_02600_),
    .S(_02841_),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_1 _08053_ (.A(_02843_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _08054_ (.A0(net3721),
    .A1(_02602_),
    .S(_02841_),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _08055_ (.A(_02844_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _08056_ (.A0(net3906),
    .A1(_02051_),
    .S(_02841_),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _08057_ (.A(_02845_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _08058_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .Y(_02846_));
 sky130_fd_sc_hd__buf_8 _08059_ (.A(_00407_),
    .X(_02847_));
 sky130_fd_sc_hd__o31a_2 _08060_ (.A1(_02846_),
    .A2(_02762_),
    .A3(_02763_),
    .B1(_02847_),
    .X(_02848_));
 sky130_fd_sc_hd__mux2_1 _08061_ (.A0(_02643_),
    .A1(net3697),
    .S(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_1 _08062_ (.A(_02849_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _08063_ (.A0(_02650_),
    .A1(net3154),
    .S(_02848_),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _08064_ (.A(_02850_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _08065_ (.A0(_02652_),
    .A1(net3922),
    .S(_02848_),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _08066_ (.A(_02851_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _08067_ (.A0(_02779_),
    .A1(net3943),
    .S(_02848_),
    .X(_02852_));
 sky130_fd_sc_hd__clkbuf_1 _08068_ (.A(_02852_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _08069_ (.A(_02762_),
    .B(_02785_),
    .X(_02853_));
 sky130_fd_sc_hd__o41a_2 _08070_ (.A1(_02772_),
    .A2(_02771_),
    .A3(_02773_),
    .A4(_02853_),
    .B1(_01497_),
    .X(_02854_));
 sky130_fd_sc_hd__mux2_1 _08071_ (.A0(_02643_),
    .A1(net3558),
    .S(_02854_),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_1 _08072_ (.A(_02855_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _08073_ (.A0(_02650_),
    .A1(net3222),
    .S(_02854_),
    .X(_02856_));
 sky130_fd_sc_hd__clkbuf_1 _08074_ (.A(_02856_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _08075_ (.A0(_02652_),
    .A1(net3311),
    .S(_02854_),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_1 _08076_ (.A(_02857_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _08077_ (.A0(_02779_),
    .A1(net3792),
    .S(_02854_),
    .X(_02858_));
 sky130_fd_sc_hd__clkbuf_1 _08078_ (.A(_02858_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _08079_ (.A(_02782_),
    .B(_02853_),
    .Y(_02859_));
 sky130_fd_sc_hd__or2_1 _08080_ (.A(net3913),
    .B(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__nand2_1 _08081_ (.A(_02787_),
    .B(_02859_),
    .Y(_02861_));
 sky130_fd_sc_hd__a31o_1 _08082_ (.A1(_02696_),
    .A2(_02860_),
    .A3(_02861_),
    .B1(_02711_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__nand2_1 _08083_ (.A(_02791_),
    .B(_02859_),
    .Y(_02862_));
 sky130_fd_sc_hd__or2_1 _08084_ (.A(net4084),
    .B(_02859_),
    .X(_02863_));
 sky130_fd_sc_hd__a31o_1 _08085_ (.A1(_02696_),
    .A2(_02862_),
    .A3(_02863_),
    .B1(_02133_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__buf_4 _08086_ (.A(_00195_),
    .X(_02864_));
 sky130_fd_sc_hd__or2_1 _08087_ (.A(net3607),
    .B(_02859_),
    .X(_02865_));
 sky130_fd_sc_hd__nand2_1 _08088_ (.A(_02794_),
    .B(_02859_),
    .Y(_02866_));
 sky130_fd_sc_hd__a31o_1 _08089_ (.A1(_02864_),
    .A2(_02865_),
    .A3(_02866_),
    .B1(_02634_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__nor2_1 _08090_ (.A(net3920),
    .B(_02859_),
    .Y(_02867_));
 sky130_fd_sc_hd__buf_6 _08091_ (.A(_00267_),
    .X(_02868_));
 sky130_fd_sc_hd__a211o_1 _08092_ (.A1(_02797_),
    .A2(_02859_),
    .B1(_02867_),
    .C1(_02868_),
    .X(_02869_));
 sky130_fd_sc_hd__nand2_1 _08093_ (.A(_02031_),
    .B(_02869_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3_2 _08094_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_02783_),
    .C(_02801_),
    .X(_02870_));
 sky130_fd_sc_hd__nor2_1 _08095_ (.A(_01971_),
    .B(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__a221o_1 _08096_ (.A1(_01762_),
    .A2(_02870_),
    .B1(_02871_),
    .B2(net3408),
    .C1(_01766_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__buf_4 _08097_ (.A(_00215_),
    .X(_02872_));
 sky130_fd_sc_hd__a221o_1 _08098_ (.A1(_01771_),
    .A2(_02870_),
    .B1(_02871_),
    .B2(net3174),
    .C1(_02872_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _08099_ (.A1(_01850_),
    .A2(_02870_),
    .B1(_02871_),
    .B2(net3211),
    .C1(_01973_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__mux4_1 _08100_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A3(_01585_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .X(_02873_));
 sky130_fd_sc_hd__mux4_1 _08101_ (.A0(_01587_),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_1 _08102_ (.A0(_02873_),
    .A1(_02874_),
    .S(net3154),
    .X(_02875_));
 sky130_fd_sc_hd__clkbuf_1 _08103_ (.A(_02875_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ));
 sky130_fd_sc_hd__mux4_1 _08104_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(_01676_),
    .A2(_01587_),
    .A3(_01588_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ),
    .X(_02876_));
 sky130_fd_sc_hd__mux4_1 _08105_ (.A0(_01678_),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _08106_ (.A0(_02876_),
    .A1(_02877_),
    .S(net3222),
    .X(_02878_));
 sky130_fd_sc_hd__clkbuf_1 _08107_ (.A(_02878_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ));
 sky130_fd_sc_hd__mux4_1 _08108_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A1(_01676_),
    .A2(_01678_),
    .A3(_01585_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .X(_02879_));
 sky130_fd_sc_hd__mux4_1 _08109_ (.A0(_01584_),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_1 _08110_ (.A0(_02879_),
    .A1(_02880_),
    .S(net3792),
    .X(_02881_));
 sky130_fd_sc_hd__clkbuf_1 _08111_ (.A(_02881_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ));
 sky130_fd_sc_hd__mux4_1 _08112_ (.A0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A3(_01585_),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ),
    .X(_02882_));
 sky130_fd_sc_hd__mux4_1 _08113_ (.A0(_01584_),
    .A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A2(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ),
    .X(_02883_));
 sky130_fd_sc_hd__mux2_1 _08114_ (.A0(_02882_),
    .A1(_02883_),
    .S(net3607),
    .X(_02884_));
 sky130_fd_sc_hd__clkbuf_1 _08115_ (.A(_02884_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ));
 sky130_fd_sc_hd__and2_1 _08116_ (.A(_01858_),
    .B(_01757_),
    .X(_02885_));
 sky130_fd_sc_hd__mux2_1 _08117_ (.A0(_02760_),
    .A1(_02885_),
    .S(_01863_),
    .X(_02886_));
 sky130_fd_sc_hd__clkbuf_1 _08118_ (.A(_02886_),
    .X(_00010_));
 sky130_fd_sc_hd__clkbuf_4 _08119_ (.A(_00171_),
    .X(_02887_));
 sky130_fd_sc_hd__nand3b_2 _08120_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .C(_01878_),
    .Y(_02888_));
 sky130_fd_sc_hd__or3_1 _08121_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_02889_));
 sky130_fd_sc_hd__or2_1 _08122_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08123_ (.A(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__o21a_1 _08124_ (.A1(_02888_),
    .A2(_02891_),
    .B1(_02092_),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_1 _08125_ (.A0(_02887_),
    .A1(net3454),
    .S(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__clkbuf_1 _08126_ (.A(_02893_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__clkbuf_4 _08127_ (.A(_00184_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _08128_ (.A0(_02894_),
    .A1(net3457),
    .S(_02892_),
    .X(_02895_));
 sky130_fd_sc_hd__clkbuf_1 _08129_ (.A(_02895_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__clkbuf_4 _08130_ (.A(_00551_),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_1 _08131_ (.A0(_02896_),
    .A1(net3524),
    .S(_02892_),
    .X(_02897_));
 sky130_fd_sc_hd__clkbuf_1 _08132_ (.A(_02897_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _08133_ (.A0(_02779_),
    .A1(net3486),
    .S(_02892_),
    .X(_02898_));
 sky130_fd_sc_hd__clkbuf_1 _08134_ (.A(_02898_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _08135_ (.A(net4165),
    .X(_02899_));
 sky130_fd_sc_hd__clkbuf_2 _08136_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .X(_02900_));
 sky130_fd_sc_hd__inv_2 _08137_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .Y(_02901_));
 sky130_fd_sc_hd__or4_1 _08138_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02900_),
    .C(_02901_),
    .D(_02888_),
    .X(_02902_));
 sky130_fd_sc_hd__o21a_1 _08139_ (.A1(_02899_),
    .A2(_02902_),
    .B1(_02092_),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_1 _08140_ (.A0(_02887_),
    .A1(net3402),
    .S(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__clkbuf_1 _08141_ (.A(_02904_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _08142_ (.A0(_02894_),
    .A1(net3545),
    .S(_02903_),
    .X(_02905_));
 sky130_fd_sc_hd__clkbuf_1 _08143_ (.A(_02905_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _08144_ (.A0(_02896_),
    .A1(net3281),
    .S(_02903_),
    .X(_02906_));
 sky130_fd_sc_hd__clkbuf_1 _08145_ (.A(_02906_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _08146_ (.A0(_02779_),
    .A1(net3368),
    .S(_02903_),
    .X(_02907_));
 sky130_fd_sc_hd__clkbuf_1 _08147_ (.A(_02907_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _08148_ (.A(_02899_),
    .Y(_02908_));
 sky130_fd_sc_hd__or3_2 _08149_ (.A(_02900_),
    .B(_02908_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_02909_));
 sky130_fd_sc_hd__and3b_1 _08150_ (.A_N(\c.genblk1.genblk1.subs.cs[2].c.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .C(_00311_),
    .X(_02910_));
 sky130_fd_sc_hd__clkbuf_2 _08151_ (.A(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__nand2_1 _08152_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02889_),
    .Y(_02912_));
 sky130_fd_sc_hd__and2_1 _08153_ (.A(_02891_),
    .B(_02912_),
    .X(_02913_));
 sky130_fd_sc_hd__nand2_1 _08154_ (.A(_02911_),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__nand2_1 _08155_ (.A(_02003_),
    .B(_02891_),
    .Y(_02915_));
 sky130_fd_sc_hd__or3_1 _08156_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02888_),
    .C(_02909_),
    .X(_02916_));
 sky130_fd_sc_hd__nand2_1 _08157_ (.A(net3346),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__o31a_1 _08158_ (.A1(_02909_),
    .A2(_02914_),
    .A3(_02915_),
    .B1(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__o21ai_1 _08159_ (.A1(_02838_),
    .A2(_02918_),
    .B1(_02145_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_1 _08160_ (.A(_00211_),
    .B(_02891_),
    .Y(_02919_));
 sky130_fd_sc_hd__nand2_1 _08161_ (.A(net3709),
    .B(_02916_),
    .Y(_02920_));
 sky130_fd_sc_hd__o31a_1 _08162_ (.A1(_02909_),
    .A2(_02914_),
    .A3(_02919_),
    .B1(_02920_),
    .X(_02921_));
 sky130_fd_sc_hd__o21ai_1 _08163_ (.A1(_02838_),
    .A2(_02921_),
    .B1(_02714_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__nand2_1 _08164_ (.A(_02573_),
    .B(_02891_),
    .Y(_02922_));
 sky130_fd_sc_hd__nand2_1 _08165_ (.A(net3634),
    .B(_02916_),
    .Y(_02923_));
 sky130_fd_sc_hd__o31a_1 _08166_ (.A1(_02909_),
    .A2(_02914_),
    .A3(_02922_),
    .B1(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__o21ai_1 _08167_ (.A1(_02838_),
    .A2(_02924_),
    .B1(_02740_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__nand2_1 _08168_ (.A(_01452_),
    .B(_02891_),
    .Y(_02925_));
 sky130_fd_sc_hd__nand2_1 _08169_ (.A(net3753),
    .B(_02916_),
    .Y(_02926_));
 sky130_fd_sc_hd__o31a_1 _08170_ (.A1(_02909_),
    .A2(_02914_),
    .A3(_02925_),
    .B1(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__buf_6 _08171_ (.A(_00226_),
    .X(_02928_));
 sky130_fd_sc_hd__o21ai_1 _08172_ (.A1(_02838_),
    .A2(_02927_),
    .B1(_02928_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_1 _08173_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_02888_),
    .Y(_02929_));
 sky130_fd_sc_hd__and3b_2 _08174_ (.A_N(_02900_),
    .B(_02899_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_02930_));
 sky130_fd_sc_hd__a21oi_2 _08175_ (.A1(_02929_),
    .A2(_02930_),
    .B1(_02686_),
    .Y(_02931_));
 sky130_fd_sc_hd__mux2_1 _08176_ (.A0(_02887_),
    .A1(net3310),
    .S(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__clkbuf_1 _08177_ (.A(_02932_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _08178_ (.A0(_02894_),
    .A1(net3349),
    .S(_02931_),
    .X(_02933_));
 sky130_fd_sc_hd__clkbuf_1 _08179_ (.A(_02933_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _08180_ (.A0(_02896_),
    .A1(net3498),
    .S(_02931_),
    .X(_02934_));
 sky130_fd_sc_hd__clkbuf_1 _08181_ (.A(_02934_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _08182_ (.A0(_02779_),
    .A1(net3333),
    .S(_02931_),
    .X(_02935_));
 sky130_fd_sc_hd__clkbuf_1 _08183_ (.A(_02935_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4_1 _08184_ (.A(_02900_),
    .B(_02908_),
    .C(_02901_),
    .D(_02929_),
    .X(_02936_));
 sky130_fd_sc_hd__clkbuf_2 _08185_ (.A(_02936_),
    .X(_02937_));
 sky130_fd_sc_hd__nand2_1 _08186_ (.A(_02915_),
    .B(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__or2_1 _08187_ (.A(net3752),
    .B(_02937_),
    .X(_02939_));
 sky130_fd_sc_hd__a31o_1 _08188_ (.A1(_02864_),
    .A2(_02938_),
    .A3(_02939_),
    .B1(_02711_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _08189_ (.A(_02919_),
    .B(_02937_),
    .Y(_02940_));
 sky130_fd_sc_hd__or2_1 _08190_ (.A(net3821),
    .B(_02937_),
    .X(_02941_));
 sky130_fd_sc_hd__a31o_1 _08191_ (.A1(_02864_),
    .A2(_02940_),
    .A3(_02941_),
    .B1(_02133_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _08192_ (.A(_02922_),
    .B(_02937_),
    .Y(_02942_));
 sky130_fd_sc_hd__or2_1 _08193_ (.A(net3376),
    .B(_02937_),
    .X(_02943_));
 sky130_fd_sc_hd__a31o_1 _08194_ (.A1(_02864_),
    .A2(_02942_),
    .A3(_02943_),
    .B1(_02634_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _08195_ (.A(net4116),
    .B(_02937_),
    .Y(_02944_));
 sky130_fd_sc_hd__a211o_1 _08196_ (.A1(_02925_),
    .A2(_02937_),
    .B1(_02944_),
    .C1(_02868_),
    .X(_02945_));
 sky130_fd_sc_hd__nand2_1 _08197_ (.A(_02031_),
    .B(_02945_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__clkbuf_8 _08198_ (.A(_00180_),
    .X(_02946_));
 sky130_fd_sc_hd__a41o_2 _08199_ (.A1(_02900_),
    .A2(_02908_),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .A4(_02929_),
    .B1(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__mux2_1 _08200_ (.A0(net4049),
    .A1(_02597_),
    .S(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__clkbuf_1 _08201_ (.A(_02948_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _08202_ (.A0(net4159),
    .A1(_02600_),
    .S(_02947_),
    .X(_02949_));
 sky130_fd_sc_hd__clkbuf_1 _08203_ (.A(_02949_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _08204_ (.A0(net3733),
    .A1(_02602_),
    .S(_02947_),
    .X(_02950_));
 sky130_fd_sc_hd__clkbuf_1 _08205_ (.A(_02950_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__buf_6 _08206_ (.A(_00191_),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_1 _08207_ (.A0(net3600),
    .A1(_02951_),
    .S(_02947_),
    .X(_02952_));
 sky130_fd_sc_hd__clkbuf_1 _08208_ (.A(_02952_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_1 _08209_ (.A(_02900_),
    .B(_02899_),
    .C(_02901_),
    .D(_02929_),
    .X(_02953_));
 sky130_fd_sc_hd__mux2_1 _08210_ (.A0(_01827_),
    .A1(_02915_),
    .S(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__o21ai_1 _08211_ (.A1(_02838_),
    .A2(_02954_),
    .B1(_02145_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _08212_ (.A0(_01830_),
    .A1(_02919_),
    .S(_02953_),
    .X(_02955_));
 sky130_fd_sc_hd__o21ai_1 _08213_ (.A1(_02838_),
    .A2(_02955_),
    .B1(_02714_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _08214_ (.A0(_01832_),
    .A1(_02922_),
    .S(_02953_),
    .X(_02956_));
 sky130_fd_sc_hd__o21ai_1 _08215_ (.A1(_02838_),
    .A2(_02956_),
    .B1(_02740_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _08216_ (.A0(_01823_),
    .A1(_02925_),
    .S(_02953_),
    .X(_02957_));
 sky130_fd_sc_hd__o21ai_1 _08217_ (.A1(_02838_),
    .A2(_02957_),
    .B1(_02928_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _08218_ (.A1(_02900_),
    .A2(_02899_),
    .A3(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .A4(_02929_),
    .B1(_02946_),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_1 _08219_ (.A0(net3790),
    .A1(_02597_),
    .S(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__clkbuf_1 _08220_ (.A(_02959_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _08221_ (.A0(net4172),
    .A1(_02600_),
    .S(_02958_),
    .X(_02960_));
 sky130_fd_sc_hd__clkbuf_1 _08222_ (.A(_02960_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _08223_ (.A0(net3637),
    .A1(_02602_),
    .S(_02958_),
    .X(_02961_));
 sky130_fd_sc_hd__clkbuf_1 _08224_ (.A(_02961_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _08225_ (.A0(net3797),
    .A1(_02951_),
    .S(_02958_),
    .X(_02962_));
 sky130_fd_sc_hd__clkbuf_1 _08226_ (.A(_02962_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _08227_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .Y(_02963_));
 sky130_fd_sc_hd__o31a_2 _08228_ (.A1(_02963_),
    .A2(_02888_),
    .A3(_02889_),
    .B1(_02847_),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_1 _08229_ (.A0(_02887_),
    .A1(net3924),
    .S(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__clkbuf_1 _08230_ (.A(_02965_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _08231_ (.A0(_02894_),
    .A1(net3197),
    .S(_02964_),
    .X(_02966_));
 sky130_fd_sc_hd__clkbuf_1 _08232_ (.A(_02966_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _08233_ (.A0(_02896_),
    .A1(net3735),
    .S(_02964_),
    .X(_02967_));
 sky130_fd_sc_hd__clkbuf_1 _08234_ (.A(_02967_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _08235_ (.A0(_02779_),
    .A1(net3635),
    .S(_02964_),
    .X(_02968_));
 sky130_fd_sc_hd__clkbuf_1 _08236_ (.A(_02968_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _08237_ (.A(_02888_),
    .B(_02913_),
    .X(_02969_));
 sky130_fd_sc_hd__o41a_2 _08238_ (.A1(_02900_),
    .A2(_02899_),
    .A3(_02901_),
    .A4(_02969_),
    .B1(_01497_),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _08239_ (.A0(_02887_),
    .A1(net3318),
    .S(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__clkbuf_1 _08240_ (.A(_02971_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _08241_ (.A0(_02894_),
    .A1(net3466),
    .S(_02970_),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_1 _08242_ (.A(_02972_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _08243_ (.A0(_02896_),
    .A1(net3643),
    .S(_02970_),
    .X(_02973_));
 sky130_fd_sc_hd__clkbuf_1 _08244_ (.A(_02973_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _08245_ (.A0(_02779_),
    .A1(net3361),
    .S(_02970_),
    .X(_02974_));
 sky130_fd_sc_hd__clkbuf_1 _08246_ (.A(_02974_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__clkbuf_4 _08247_ (.A(_01764_),
    .X(_02975_));
 sky130_fd_sc_hd__nor2_2 _08248_ (.A(_02909_),
    .B(_02969_),
    .Y(_02976_));
 sky130_fd_sc_hd__mux2_1 _08249_ (.A0(_02751_),
    .A1(_02915_),
    .S(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__buf_6 _08250_ (.A(_00237_),
    .X(_02978_));
 sky130_fd_sc_hd__o21ai_1 _08251_ (.A1(_02975_),
    .A2(_02977_),
    .B1(_02978_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__nand2_1 _08252_ (.A(_02919_),
    .B(_02976_),
    .Y(_02979_));
 sky130_fd_sc_hd__or2_1 _08253_ (.A(net4119),
    .B(_02976_),
    .X(_02980_));
 sky130_fd_sc_hd__a31o_1 _08254_ (.A1(_02864_),
    .A2(_02979_),
    .A3(_02980_),
    .B1(_02133_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__nand2_1 _08255_ (.A(_02922_),
    .B(_02976_),
    .Y(_02981_));
 sky130_fd_sc_hd__or2_1 _08256_ (.A(net3394),
    .B(_02976_),
    .X(_02982_));
 sky130_fd_sc_hd__a31o_1 _08257_ (.A1(_02864_),
    .A2(_02981_),
    .A3(_02982_),
    .B1(_02634_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__mux2_1 _08258_ (.A0(_02755_),
    .A1(_02925_),
    .S(_02976_),
    .X(_02983_));
 sky130_fd_sc_hd__o21ai_1 _08259_ (.A1(_02975_),
    .A2(_02983_),
    .B1(_02928_),
    .Y(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3b_1 _08260_ (.A_N(_02913_),
    .B(_02930_),
    .C(_02911_),
    .X(_02984_));
 sky130_fd_sc_hd__a31oi_4 _08261_ (.A1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .A2(_02911_),
    .A3(_02930_),
    .B1(_02637_),
    .Y(_02985_));
 sky130_fd_sc_hd__a221o_1 _08262_ (.A1(_01762_),
    .A2(_02984_),
    .B1(_02985_),
    .B2(net3535),
    .C1(_00209_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _08263_ (.A1(_01771_),
    .A2(_02984_),
    .B1(_02985_),
    .B2(net3242),
    .C1(_02872_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _08264_ (.A1(_01850_),
    .A2(_02984_),
    .B1(_02985_),
    .B2(net3186),
    .C1(_01973_),
    .X(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__mux4_1 _08265_ (.A0(_00879_),
    .A1(_00881_),
    .A2(_00882_),
    .A3(_00883_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .X(_02986_));
 sky130_fd_sc_hd__clkinv_2 _08266_ (.A(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__mux4_1 _08267_ (.A0(_00886_),
    .A1(_00887_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _08268_ (.A0(_02987_),
    .A1(_02988_),
    .S(net3202),
    .X(_02989_));
 sky130_fd_sc_hd__clkbuf_1 _08269_ (.A(_02989_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ));
 sky130_fd_sc_hd__mux4_1 _08270_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(_00973_),
    .A2(_00886_),
    .A3(_00887_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(_02990_));
 sky130_fd_sc_hd__mux4_1 _08271_ (.A0(_00975_),
    .A1(_00976_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_1 _08272_ (.A0(_02990_),
    .A1(_02991_),
    .S(net3625),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_1 _08273_ (.A(_02992_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ));
 sky130_fd_sc_hd__mux4_1 _08274_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A1(_00973_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A3(_00976_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ),
    .X(_02993_));
 sky130_fd_sc_hd__mux4_1 _08275_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(_00887_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_1 _08276_ (.A0(_02993_),
    .A1(_02994_),
    .S(net3386),
    .X(_02995_));
 sky130_fd_sc_hd__clkbuf_1 _08277_ (.A(_02995_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ));
 sky130_fd_sc_hd__mux4_1 _08278_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A3(_00976_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .S1(net3804),
    .X(_02996_));
 sky130_fd_sc_hd__mux4_1 _08279_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .S1(net3804),
    .X(_02997_));
 sky130_fd_sc_hd__mux2_1 _08280_ (.A0(_02996_),
    .A1(_02997_),
    .S(net3520),
    .X(_02998_));
 sky130_fd_sc_hd__clkbuf_1 _08281_ (.A(_02998_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ));
 sky130_fd_sc_hd__mux2_1 _08282_ (.A0(_02640_),
    .A1(_02885_),
    .S(_02525_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_1 _08283_ (.A(_02999_),
    .X(_00011_));
 sky130_fd_sc_hd__nand3b_2 _08284_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .B(_01415_),
    .C(\c.genblk1.genblk1.subs.c0.cfgd ),
    .Y(_03000_));
 sky130_fd_sc_hd__or3_1 _08285_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_03001_));
 sky130_fd_sc_hd__or2_1 _08286_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08287_ (.A(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__o21a_2 _08288_ (.A1(_03000_),
    .A2(_03003_),
    .B1(_02092_),
    .X(_03004_));
 sky130_fd_sc_hd__mux2_1 _08289_ (.A0(_02887_),
    .A1(net3549),
    .S(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__clkbuf_1 _08290_ (.A(_03005_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _08291_ (.A0(_02894_),
    .A1(net3465),
    .S(_03004_),
    .X(_03006_));
 sky130_fd_sc_hd__clkbuf_1 _08292_ (.A(_03006_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _08293_ (.A0(_02896_),
    .A1(net3334),
    .S(_03004_),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_1 _08294_ (.A(_03007_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _08295_ (.A0(_02779_),
    .A1(net3409),
    .S(_03004_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_1 _08296_ (.A(_03008_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _08297_ (.A(net4150),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_2 _08298_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ),
    .X(_03010_));
 sky130_fd_sc_hd__inv_2 _08299_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .Y(_03011_));
 sky130_fd_sc_hd__or4_1 _08300_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_03010_),
    .C(_03011_),
    .D(_03000_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_8 _08301_ (.A(_00407_),
    .X(_03013_));
 sky130_fd_sc_hd__o21a_2 _08302_ (.A1(_03009_),
    .A2(_03012_),
    .B1(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_1 _08303_ (.A0(_02887_),
    .A1(net3238),
    .S(_03014_),
    .X(_03015_));
 sky130_fd_sc_hd__clkbuf_1 _08304_ (.A(_03015_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _08305_ (.A0(_02894_),
    .A1(net3150),
    .S(_03014_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_1 _08306_ (.A(_03016_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _08307_ (.A0(_02896_),
    .A1(net3151),
    .S(_03014_),
    .X(_03017_));
 sky130_fd_sc_hd__clkbuf_1 _08308_ (.A(_03017_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__clkbuf_4 _08309_ (.A(_00191_),
    .X(_03018_));
 sky130_fd_sc_hd__mux2_1 _08310_ (.A0(_03018_),
    .A1(net3525),
    .S(_03014_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_1 _08311_ (.A(_03019_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _08312_ (.A(_03009_),
    .Y(_03020_));
 sky130_fd_sc_hd__or3_1 _08313_ (.A(_03010_),
    .B(_03020_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_03021_));
 sky130_fd_sc_hd__and3b_2 _08314_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .B(_00311_),
    .C(\c.genblk1.genblk1.subs.c0.cfgd ),
    .X(_03022_));
 sky130_fd_sc_hd__nand2_1 _08315_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_03001_),
    .Y(_03023_));
 sky130_fd_sc_hd__and2_1 _08316_ (.A(_03003_),
    .B(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__nand2_1 _08317_ (.A(_03022_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__nand2_1 _08318_ (.A(_02003_),
    .B(_03003_),
    .Y(_03026_));
 sky130_fd_sc_hd__or3_1 _08319_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_03000_),
    .C(_03021_),
    .X(_03027_));
 sky130_fd_sc_hd__nand2_1 _08320_ (.A(net3710),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__o31a_1 _08321_ (.A1(_03021_),
    .A2(_03025_),
    .A3(_03026_),
    .B1(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__o21ai_1 _08322_ (.A1(_02975_),
    .A2(_03029_),
    .B1(_02978_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_1 _08323_ (.A(_01446_),
    .B(_03003_),
    .Y(_03030_));
 sky130_fd_sc_hd__or2_1 _08324_ (.A(_03021_),
    .B(_03025_),
    .X(_03031_));
 sky130_fd_sc_hd__a2bb2o_1 _08325_ (.A1_N(_03030_),
    .A2_N(_03031_),
    .B1(net3895),
    .B2(_03027_),
    .X(_03032_));
 sky130_fd_sc_hd__a21o_1 _08326_ (.A1(_02044_),
    .A2(_03032_),
    .B1(_00216_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__nand2_1 _08327_ (.A(_02573_),
    .B(_03003_),
    .Y(_03033_));
 sky130_fd_sc_hd__a2bb2o_1 _08328_ (.A1_N(_03031_),
    .A2_N(_03033_),
    .B1(net3762),
    .B2(_03027_),
    .X(_03034_));
 sky130_fd_sc_hd__a21o_1 _08329_ (.A1(_02044_),
    .A2(_03034_),
    .B1(_00262_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__nand2_1 _08330_ (.A(_01452_),
    .B(_03003_),
    .Y(_03035_));
 sky130_fd_sc_hd__o2bb2a_1 _08331_ (.A1_N(net4058),
    .A2_N(_03027_),
    .B1(_03031_),
    .B2(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__o21ai_1 _08332_ (.A1(_02975_),
    .A2(_03036_),
    .B1(_02928_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _08333_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_03000_),
    .Y(_03037_));
 sky130_fd_sc_hd__and3b_2 _08334_ (.A_N(_03010_),
    .B(_03009_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_03038_));
 sky130_fd_sc_hd__a21oi_4 _08335_ (.A1(_03037_),
    .A2(_03038_),
    .B1(_02686_),
    .Y(_03039_));
 sky130_fd_sc_hd__mux2_1 _08336_ (.A0(_02887_),
    .A1(net3369),
    .S(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__clkbuf_1 _08337_ (.A(_03040_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _08338_ (.A0(_02894_),
    .A1(net3356),
    .S(_03039_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_1 _08339_ (.A(_03041_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _08340_ (.A0(_02896_),
    .A1(net3397),
    .S(_03039_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _08341_ (.A(_03042_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _08342_ (.A0(_03018_),
    .A1(net3543),
    .S(_03039_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _08343_ (.A(_03043_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4_1 _08344_ (.A(_03010_),
    .B(_03020_),
    .C(_03011_),
    .D(_03037_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_2 _08345_ (.A(_03044_),
    .X(_03045_));
 sky130_fd_sc_hd__nand2_1 _08346_ (.A(_03026_),
    .B(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__or2_1 _08347_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .B(_03045_),
    .X(_03047_));
 sky130_fd_sc_hd__a31o_1 _08348_ (.A1(_02864_),
    .A2(_03046_),
    .A3(_03047_),
    .B1(_02711_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _08349_ (.A(_03030_),
    .B(_03045_),
    .Y(_03048_));
 sky130_fd_sc_hd__or2_1 _08350_ (.A(net4162),
    .B(_03045_),
    .X(_03049_));
 sky130_fd_sc_hd__buf_6 _08351_ (.A(_00215_),
    .X(_03050_));
 sky130_fd_sc_hd__a31o_1 _08352_ (.A1(_02864_),
    .A2(_03048_),
    .A3(_03049_),
    .B1(_03050_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _08353_ (.A(_03033_),
    .B(_03045_),
    .Y(_03051_));
 sky130_fd_sc_hd__or2_1 _08354_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .B(_03045_),
    .X(_03052_));
 sky130_fd_sc_hd__a31o_1 _08355_ (.A1(_02864_),
    .A2(_03051_),
    .A3(_03052_),
    .B1(_02634_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _08356_ (.A(net3492),
    .B(_03045_),
    .Y(_03053_));
 sky130_fd_sc_hd__a211o_1 _08357_ (.A1(_03035_),
    .A2(_03045_),
    .B1(_03053_),
    .C1(_02868_),
    .X(_03054_));
 sky130_fd_sc_hd__nand2_1 _08358_ (.A(_02031_),
    .B(_03054_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _08359_ (.A1(_03010_),
    .A2(_03020_),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .A4(_03037_),
    .B1(_02946_),
    .X(_03055_));
 sky130_fd_sc_hd__mux2_1 _08360_ (.A0(net3959),
    .A1(_02597_),
    .S(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__clkbuf_1 _08361_ (.A(_03056_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _08362_ (.A0(net4141),
    .A1(_02600_),
    .S(_03055_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_1 _08363_ (.A(_03057_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _08364_ (.A0(net3908),
    .A1(_02602_),
    .S(_03055_),
    .X(_03058_));
 sky130_fd_sc_hd__clkbuf_1 _08365_ (.A(_03058_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _08366_ (.A0(net3813),
    .A1(_02951_),
    .S(_03055_),
    .X(_03059_));
 sky130_fd_sc_hd__clkbuf_1 _08367_ (.A(_03059_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_1 _08368_ (.A(_03010_),
    .B(_03009_),
    .C(_03011_),
    .D(_03037_),
    .X(_03060_));
 sky130_fd_sc_hd__or2_1 _08369_ (.A(net4192),
    .B(_03060_),
    .X(_03061_));
 sky130_fd_sc_hd__nand2_1 _08370_ (.A(_03026_),
    .B(_03060_),
    .Y(_03062_));
 sky130_fd_sc_hd__a31o_1 _08371_ (.A1(_02864_),
    .A2(_03061_),
    .A3(_03062_),
    .B1(_02711_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _08372_ (.A0(_02157_),
    .A1(_03030_),
    .S(_03060_),
    .X(_03063_));
 sky130_fd_sc_hd__o21ai_1 _08373_ (.A1(_02975_),
    .A2(_03063_),
    .B1(_02714_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _08374_ (.A0(_02159_),
    .A1(_03033_),
    .S(_03060_),
    .X(_03064_));
 sky130_fd_sc_hd__o21ai_1 _08375_ (.A1(_02975_),
    .A2(_03064_),
    .B1(_02740_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _08376_ (.A0(_02165_),
    .A1(_03035_),
    .S(_03060_),
    .X(_03065_));
 sky130_fd_sc_hd__o21ai_1 _08377_ (.A1(_02975_),
    .A2(_03065_),
    .B1(_02928_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _08378_ (.A1(_03010_),
    .A2(_03009_),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .A4(_03037_),
    .B1(_02946_),
    .X(_03066_));
 sky130_fd_sc_hd__mux2_1 _08379_ (.A0(net4115),
    .A1(_02597_),
    .S(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__clkbuf_1 _08380_ (.A(_03067_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _08381_ (.A0(net3903),
    .A1(_02600_),
    .S(_03066_),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_1 _08382_ (.A(_03068_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _08383_ (.A0(net3583),
    .A1(_02602_),
    .S(_03066_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _08384_ (.A(_03069_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _08385_ (.A0(net4020),
    .A1(_02951_),
    .S(_03066_),
    .X(_03070_));
 sky130_fd_sc_hd__clkbuf_1 _08386_ (.A(_03070_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _08387_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .Y(_03071_));
 sky130_fd_sc_hd__o31a_2 _08388_ (.A1(_03071_),
    .A2(_03000_),
    .A3(_03001_),
    .B1(_02847_),
    .X(_03072_));
 sky130_fd_sc_hd__mux2_1 _08389_ (.A0(_02887_),
    .A1(net3758),
    .S(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_1 _08390_ (.A(_03073_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _08391_ (.A0(_02894_),
    .A1(net3291),
    .S(_03072_),
    .X(_03074_));
 sky130_fd_sc_hd__clkbuf_1 _08392_ (.A(_03074_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _08393_ (.A0(_02896_),
    .A1(net3597),
    .S(_03072_),
    .X(_03075_));
 sky130_fd_sc_hd__clkbuf_1 _08394_ (.A(_03075_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _08395_ (.A0(_03018_),
    .A1(net3996),
    .S(_03072_),
    .X(_03076_));
 sky130_fd_sc_hd__clkbuf_1 _08396_ (.A(_03076_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _08397_ (.A(_03000_),
    .B(_03024_),
    .X(_03077_));
 sky130_fd_sc_hd__o41a_2 _08398_ (.A1(_03010_),
    .A2(_03009_),
    .A3(_03011_),
    .A4(_03077_),
    .B1(_01497_),
    .X(_03078_));
 sky130_fd_sc_hd__mux2_1 _08399_ (.A0(_02887_),
    .A1(net3881),
    .S(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__clkbuf_1 _08400_ (.A(_03079_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _08401_ (.A0(_02894_),
    .A1(net3331),
    .S(_03078_),
    .X(_03080_));
 sky130_fd_sc_hd__clkbuf_1 _08402_ (.A(_03080_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _08403_ (.A0(_02896_),
    .A1(net3910),
    .S(_03078_),
    .X(_03081_));
 sky130_fd_sc_hd__clkbuf_1 _08404_ (.A(_03081_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _08405_ (.A0(_03018_),
    .A1(net3681),
    .S(_03078_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_1 _08406_ (.A(_03082_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _08407_ (.A(_03021_),
    .B(_03077_),
    .Y(_03083_));
 sky130_fd_sc_hd__mux2_1 _08408_ (.A0(_02540_),
    .A1(_03026_),
    .S(_03083_),
    .X(_03084_));
 sky130_fd_sc_hd__o21ai_1 _08409_ (.A1(_02975_),
    .A2(_03084_),
    .B1(_02978_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__buf_4 _08410_ (.A(_00195_),
    .X(_03085_));
 sky130_fd_sc_hd__nand2_1 _08411_ (.A(_03030_),
    .B(_03083_),
    .Y(_03086_));
 sky130_fd_sc_hd__or2_1 _08412_ (.A(net4000),
    .B(_03083_),
    .X(_03087_));
 sky130_fd_sc_hd__a31o_1 _08413_ (.A1(_03085_),
    .A2(_03086_),
    .A3(_03087_),
    .B1(_03050_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__or2_1 _08414_ (.A(net3223),
    .B(_03083_),
    .X(_03088_));
 sky130_fd_sc_hd__nand2_1 _08415_ (.A(_03033_),
    .B(_03083_),
    .Y(_03089_));
 sky130_fd_sc_hd__a31o_1 _08416_ (.A1(_03085_),
    .A2(_03088_),
    .A3(_03089_),
    .B1(_02634_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__mux2_1 _08417_ (.A0(_02546_),
    .A1(_03035_),
    .S(_03083_),
    .X(_03090_));
 sky130_fd_sc_hd__o21ai_1 _08418_ (.A1(_02975_),
    .A2(_03090_),
    .B1(_02928_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3b_1 _08419_ (.A_N(_03024_),
    .B(_03038_),
    .C(_03022_),
    .X(_03091_));
 sky130_fd_sc_hd__a31oi_4 _08420_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .A2(_03022_),
    .A3(_03038_),
    .B1(_02637_),
    .Y(_03092_));
 sky130_fd_sc_hd__a221o_1 _08421_ (.A1(_01762_),
    .A2(_03091_),
    .B1(_03092_),
    .B2(net3243),
    .C1(_00209_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _08422_ (.A1(_01771_),
    .A2(_03091_),
    .B1(_03092_),
    .B2(net3213),
    .C1(_02872_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _08423_ (.A1(_01850_),
    .A2(_03091_),
    .B1(_03092_),
    .B2(net3305),
    .C1(_01973_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__mux4_1 _08424_ (.A0(_00879_),
    .A1(_00881_),
    .A2(_00882_),
    .A3(_00883_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .X(_03093_));
 sky130_fd_sc_hd__clkinv_2 _08425_ (.A(_03093_),
    .Y(_03094_));
 sky130_fd_sc_hd__mux4_1 _08426_ (.A0(_00886_),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .X(_03095_));
 sky130_fd_sc_hd__mux2_1 _08427_ (.A0(_03094_),
    .A1(_03095_),
    .S(net3195),
    .X(_03096_));
 sky130_fd_sc_hd__clkbuf_1 _08428_ (.A(_03096_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ));
 sky130_fd_sc_hd__mux4_1 _08429_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ),
    .A2(_00886_),
    .A3(_00887_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(_03097_));
 sky130_fd_sc_hd__mux4_1 _08430_ (.A0(_00975_),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(_03098_));
 sky130_fd_sc_hd__mux2_1 _08431_ (.A0(net3373),
    .A1(_03098_),
    .S(net3321),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_1 _08432_ (.A(_03099_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ));
 sky130_fd_sc_hd__mux4_1 _08433_ (.A0(_00975_),
    .A1(_00976_),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A3(_00973_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .S1(_01961_),
    .X(_03100_));
 sky130_fd_sc_hd__mux4_1 _08434_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A3(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .X(_03101_));
 sky130_fd_sc_hd__mux2_1 _08435_ (.A0(_03100_),
    .A1(_03101_),
    .S(net3682),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_1 _08436_ (.A(_03102_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ));
 sky130_fd_sc_hd__and2_2 _08437_ (.A(_01858_),
    .B(_02489_),
    .X(_03103_));
 sky130_fd_sc_hd__and2_1 _08438_ (.A(_01578_),
    .B(_02224_),
    .X(_03104_));
 sky130_fd_sc_hd__mux2_1 _08439_ (.A0(_03103_),
    .A1(_03104_),
    .S(_01863_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_1 _08440_ (.A(_03105_),
    .X(_00004_));
 sky130_fd_sc_hd__mux4_1 _08441_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(_00886_),
    .A2(_00888_),
    .A3(_00889_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .S1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .X(_03106_));
 sky130_fd_sc_hd__mux4_1 _08442_ (.A0(_00975_),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A3(_00973_),
    .S0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .S1(_01968_),
    .X(_03107_));
 sky130_fd_sc_hd__mux2_1 _08443_ (.A0(_03106_),
    .A1(_03107_),
    .S(_01966_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _08444_ (.A(_03108_),
    .X(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ));
 sky130_fd_sc_hd__clkbuf_4 _08445_ (.A(_00171_),
    .X(_03109_));
 sky130_fd_sc_hd__nand3b_2 _08446_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .C(_01878_),
    .Y(_03110_));
 sky130_fd_sc_hd__or3_1 _08447_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_03111_));
 sky130_fd_sc_hd__or2_1 _08448_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03111_),
    .X(_03112_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08449_ (.A(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__o21a_2 _08450_ (.A1(_03110_),
    .A2(_03113_),
    .B1(_03013_),
    .X(_03114_));
 sky130_fd_sc_hd__mux2_1 _08451_ (.A0(_03109_),
    .A1(net3737),
    .S(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__clkbuf_1 _08452_ (.A(_03115_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__clkbuf_4 _08453_ (.A(_00184_),
    .X(_03116_));
 sky130_fd_sc_hd__mux2_1 _08454_ (.A0(_03116_),
    .A1(net3666),
    .S(_03114_),
    .X(_03117_));
 sky130_fd_sc_hd__clkbuf_1 _08455_ (.A(_03117_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__buf_4 _08456_ (.A(_00551_),
    .X(_03118_));
 sky130_fd_sc_hd__mux2_1 _08457_ (.A0(_03118_),
    .A1(net3537),
    .S(_03114_),
    .X(_03119_));
 sky130_fd_sc_hd__clkbuf_1 _08458_ (.A(_03119_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _08459_ (.A0(_03018_),
    .A1(net3503),
    .S(_03114_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_1 _08460_ (.A(_03120_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _08461_ (.A(net4169),
    .X(_03121_));
 sky130_fd_sc_hd__clkbuf_2 _08462_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ),
    .X(_03122_));
 sky130_fd_sc_hd__inv_2 _08463_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .Y(_03123_));
 sky130_fd_sc_hd__or4_1 _08464_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03122_),
    .C(_03123_),
    .D(_03110_),
    .X(_03124_));
 sky130_fd_sc_hd__o21a_1 _08465_ (.A1(_03121_),
    .A2(_03124_),
    .B1(_03013_),
    .X(_03125_));
 sky130_fd_sc_hd__mux2_1 _08466_ (.A0(_03109_),
    .A1(net3611),
    .S(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__clkbuf_1 _08467_ (.A(_03126_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _08468_ (.A0(_03116_),
    .A1(net3159),
    .S(_03125_),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_1 _08469_ (.A(_03127_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _08470_ (.A0(_03118_),
    .A1(net3273),
    .S(_03125_),
    .X(_03128_));
 sky130_fd_sc_hd__clkbuf_1 _08471_ (.A(_03128_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _08472_ (.A0(_03018_),
    .A1(net3352),
    .S(_03125_),
    .X(_03129_));
 sky130_fd_sc_hd__clkbuf_1 _08473_ (.A(_03129_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _08474_ (.A(_03121_),
    .Y(_03130_));
 sky130_fd_sc_hd__or3_2 _08475_ (.A(_03122_),
    .B(_03130_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_03131_));
 sky130_fd_sc_hd__and3b_1 _08476_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .C(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ),
    .X(_03132_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08477_ (.A(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__nand2_1 _08478_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03111_),
    .Y(_03134_));
 sky130_fd_sc_hd__and2_1 _08479_ (.A(_03113_),
    .B(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__nand2_1 _08480_ (.A(_03133_),
    .B(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__nand2_1 _08481_ (.A(_02003_),
    .B(_03113_),
    .Y(_03137_));
 sky130_fd_sc_hd__or3_1 _08482_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03110_),
    .C(_03131_),
    .X(_03138_));
 sky130_fd_sc_hd__nand2_1 _08483_ (.A(net3703),
    .B(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__o31a_1 _08484_ (.A1(_03131_),
    .A2(_03136_),
    .A3(_03137_),
    .B1(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__o21ai_1 _08485_ (.A1(_02975_),
    .A2(_03140_),
    .B1(_02978_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__buf_2 _08486_ (.A(_01764_),
    .X(_03141_));
 sky130_fd_sc_hd__nand2_1 _08487_ (.A(_00211_),
    .B(_03113_),
    .Y(_03142_));
 sky130_fd_sc_hd__nand2_1 _08488_ (.A(net3675),
    .B(_03138_),
    .Y(_03143_));
 sky130_fd_sc_hd__o31a_1 _08489_ (.A1(_03131_),
    .A2(_03136_),
    .A3(_03142_),
    .B1(_03143_),
    .X(_03144_));
 sky130_fd_sc_hd__o21ai_1 _08490_ (.A1(_03141_),
    .A2(_03144_),
    .B1(_02714_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__nand2_1 _08491_ (.A(_02573_),
    .B(_03113_),
    .Y(_03145_));
 sky130_fd_sc_hd__nand2_1 _08492_ (.A(net3741),
    .B(_03138_),
    .Y(_03146_));
 sky130_fd_sc_hd__o31a_1 _08493_ (.A1(_03131_),
    .A2(_03136_),
    .A3(_03145_),
    .B1(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__o21ai_1 _08494_ (.A1(_03141_),
    .A2(_03147_),
    .B1(_02740_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__nand2_1 _08495_ (.A(_00264_),
    .B(_03113_),
    .Y(_03148_));
 sky130_fd_sc_hd__nand2_1 _08496_ (.A(net3699),
    .B(_03138_),
    .Y(_03149_));
 sky130_fd_sc_hd__o31a_1 _08497_ (.A1(_03131_),
    .A2(_03136_),
    .A3(_03148_),
    .B1(_03149_),
    .X(_03150_));
 sky130_fd_sc_hd__o21ai_1 _08498_ (.A1(_03141_),
    .A2(_03150_),
    .B1(_02928_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_1 _08499_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03110_),
    .Y(_03151_));
 sky130_fd_sc_hd__and3b_1 _08500_ (.A_N(_03122_),
    .B(_03121_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_03152_));
 sky130_fd_sc_hd__a21oi_2 _08501_ (.A1(_03151_),
    .A2(_03152_),
    .B1(_02686_),
    .Y(_03153_));
 sky130_fd_sc_hd__mux2_1 _08502_ (.A0(_03109_),
    .A1(net3363),
    .S(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__clkbuf_1 _08503_ (.A(_03154_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _08504_ (.A0(_03116_),
    .A1(net3451),
    .S(_03153_),
    .X(_03155_));
 sky130_fd_sc_hd__clkbuf_1 _08505_ (.A(_03155_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _08506_ (.A0(_03118_),
    .A1(net3328),
    .S(_03153_),
    .X(_03156_));
 sky130_fd_sc_hd__clkbuf_1 _08507_ (.A(_03156_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _08508_ (.A0(_03018_),
    .A1(net3656),
    .S(_03153_),
    .X(_03157_));
 sky130_fd_sc_hd__clkbuf_1 _08509_ (.A(_03157_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4_1 _08510_ (.A(_03122_),
    .B(_03130_),
    .C(_03123_),
    .D(_03151_),
    .X(_03158_));
 sky130_fd_sc_hd__clkbuf_2 _08511_ (.A(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__nand2_1 _08512_ (.A(_03137_),
    .B(_03159_),
    .Y(_03160_));
 sky130_fd_sc_hd__or2_1 _08513_ (.A(net3883),
    .B(_03159_),
    .X(_03161_));
 sky130_fd_sc_hd__a31o_1 _08514_ (.A1(_03085_),
    .A2(_03160_),
    .A3(_03161_),
    .B1(_02711_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _08515_ (.A(_03142_),
    .B(_03159_),
    .Y(_03162_));
 sky130_fd_sc_hd__or2_1 _08516_ (.A(net3989),
    .B(_03159_),
    .X(_03163_));
 sky130_fd_sc_hd__a31o_1 _08517_ (.A1(_03085_),
    .A2(_03162_),
    .A3(_03163_),
    .B1(_03050_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _08518_ (.A(_03145_),
    .B(_03159_),
    .Y(_03164_));
 sky130_fd_sc_hd__or2_1 _08519_ (.A(net3297),
    .B(_03159_),
    .X(_03165_));
 sky130_fd_sc_hd__a31o_1 _08520_ (.A1(_03085_),
    .A2(_03164_),
    .A3(_03165_),
    .B1(_02634_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__buf_6 _08521_ (.A(_00227_),
    .X(_03166_));
 sky130_fd_sc_hd__nor2_1 _08522_ (.A(net3954),
    .B(_03159_),
    .Y(_03167_));
 sky130_fd_sc_hd__a211o_1 _08523_ (.A1(_03148_),
    .A2(_03159_),
    .B1(_03167_),
    .C1(_02868_),
    .X(_03168_));
 sky130_fd_sc_hd__nand2_1 _08524_ (.A(_03166_),
    .B(_03168_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__buf_4 _08525_ (.A(_00235_),
    .X(_03169_));
 sky130_fd_sc_hd__a41o_2 _08526_ (.A1(_03122_),
    .A2(_03130_),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .A4(_03151_),
    .B1(_02946_),
    .X(_03170_));
 sky130_fd_sc_hd__mux2_1 _08527_ (.A0(net4088),
    .A1(_03169_),
    .S(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__clkbuf_1 _08528_ (.A(_03171_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__clkbuf_8 _08529_ (.A(_00292_),
    .X(_03172_));
 sky130_fd_sc_hd__mux2_1 _08530_ (.A0(net3962),
    .A1(_03172_),
    .S(_03170_),
    .X(_03173_));
 sky130_fd_sc_hd__clkbuf_1 _08531_ (.A(_03173_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__buf_4 _08532_ (.A(_00188_),
    .X(_03174_));
 sky130_fd_sc_hd__mux2_1 _08533_ (.A0(net3685),
    .A1(_03174_),
    .S(_03170_),
    .X(_03175_));
 sky130_fd_sc_hd__clkbuf_1 _08534_ (.A(_03175_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _08535_ (.A0(net3210),
    .A1(_02951_),
    .S(_03170_),
    .X(_03176_));
 sky130_fd_sc_hd__clkbuf_1 _08536_ (.A(_03176_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_1 _08537_ (.A(_03122_),
    .B(_03121_),
    .C(_03123_),
    .D(_03151_),
    .X(_03177_));
 sky130_fd_sc_hd__mux2_1 _08538_ (.A0(_02265_),
    .A1(_03137_),
    .S(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__o21ai_1 _08539_ (.A1(_03141_),
    .A2(_03178_),
    .B1(_02978_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _08540_ (.A0(_02268_),
    .A1(_03142_),
    .S(_03177_),
    .X(_03179_));
 sky130_fd_sc_hd__o21ai_1 _08541_ (.A1(_03141_),
    .A2(_03179_),
    .B1(_02714_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _08542_ (.A0(_02263_),
    .A1(_03145_),
    .S(_03177_),
    .X(_03180_));
 sky130_fd_sc_hd__o21ai_1 _08543_ (.A1(_03141_),
    .A2(_03180_),
    .B1(_02740_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _08544_ (.A0(_02260_),
    .A1(_03148_),
    .S(_03177_),
    .X(_03181_));
 sky130_fd_sc_hd__o21ai_1 _08545_ (.A1(_03141_),
    .A2(_03181_),
    .B1(_02928_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _08546_ (.A1(_03122_),
    .A2(_03121_),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .A4(_03151_),
    .B1(_02946_),
    .X(_03182_));
 sky130_fd_sc_hd__mux2_1 _08547_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .A1(_03169_),
    .S(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__clkbuf_1 _08548_ (.A(_03183_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _08549_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A1(_03172_),
    .S(_03182_),
    .X(_03184_));
 sky130_fd_sc_hd__clkbuf_1 _08550_ (.A(_03184_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _08551_ (.A0(net3653),
    .A1(_03174_),
    .S(_03182_),
    .X(_03185_));
 sky130_fd_sc_hd__clkbuf_1 _08552_ (.A(_03185_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _08553_ (.A0(net3965),
    .A1(_02951_),
    .S(_03182_),
    .X(_03186_));
 sky130_fd_sc_hd__clkbuf_1 _08554_ (.A(_03186_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _08555_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .Y(_03187_));
 sky130_fd_sc_hd__o31a_2 _08556_ (.A1(_03187_),
    .A2(_03110_),
    .A3(_03111_),
    .B1(_02847_),
    .X(_03188_));
 sky130_fd_sc_hd__mux2_1 _08557_ (.A0(_03109_),
    .A1(net3638),
    .S(_03188_),
    .X(_03189_));
 sky130_fd_sc_hd__clkbuf_1 _08558_ (.A(_03189_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _08559_ (.A0(_03116_),
    .A1(net3365),
    .S(_03188_),
    .X(_03190_));
 sky130_fd_sc_hd__clkbuf_1 _08560_ (.A(_03190_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _08561_ (.A0(_03118_),
    .A1(net3921),
    .S(_03188_),
    .X(_03191_));
 sky130_fd_sc_hd__clkbuf_1 _08562_ (.A(_03191_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _08563_ (.A0(_03018_),
    .A1(net3969),
    .S(_03188_),
    .X(_03192_));
 sky130_fd_sc_hd__clkbuf_1 _08564_ (.A(_03192_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _08565_ (.A(_03110_),
    .B(_03135_),
    .X(_03193_));
 sky130_fd_sc_hd__o41a_2 _08566_ (.A1(_03122_),
    .A2(_03121_),
    .A3(_03123_),
    .A4(_03193_),
    .B1(_01497_),
    .X(_03194_));
 sky130_fd_sc_hd__mux2_1 _08567_ (.A0(_03109_),
    .A1(net3911),
    .S(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__clkbuf_1 _08568_ (.A(_03195_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _08569_ (.A0(_03116_),
    .A1(net3232),
    .S(_03194_),
    .X(_03196_));
 sky130_fd_sc_hd__clkbuf_1 _08570_ (.A(_03196_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _08571_ (.A0(_03118_),
    .A1(net3290),
    .S(_03194_),
    .X(_03197_));
 sky130_fd_sc_hd__clkbuf_1 _08572_ (.A(_03197_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _08573_ (.A0(_03018_),
    .A1(net3156),
    .S(_03194_),
    .X(_03198_));
 sky130_fd_sc_hd__clkbuf_1 _08574_ (.A(_03198_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _08575_ (.A(_03131_),
    .B(_03193_),
    .Y(_03199_));
 sky130_fd_sc_hd__or2_1 _08576_ (.A(net3950),
    .B(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__nand2_1 _08577_ (.A(_03137_),
    .B(_03199_),
    .Y(_03201_));
 sky130_fd_sc_hd__a31o_1 _08578_ (.A1(_03085_),
    .A2(_03200_),
    .A3(_03201_),
    .B1(_02711_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__nand2_1 _08579_ (.A(_03142_),
    .B(_03199_),
    .Y(_03202_));
 sky130_fd_sc_hd__or2_1 _08580_ (.A(net3961),
    .B(_03199_),
    .X(_03203_));
 sky130_fd_sc_hd__a31o_1 _08581_ (.A1(_03085_),
    .A2(_03202_),
    .A3(_03203_),
    .B1(_03050_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__or2_1 _08582_ (.A(net3585),
    .B(_03199_),
    .X(_03204_));
 sky130_fd_sc_hd__nand2_1 _08583_ (.A(_03145_),
    .B(_03199_),
    .Y(_03205_));
 sky130_fd_sc_hd__a31o_1 _08584_ (.A1(_03085_),
    .A2(_03204_),
    .A3(_03205_),
    .B1(_02634_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__nor2_1 _08585_ (.A(net4033),
    .B(_03199_),
    .Y(_03206_));
 sky130_fd_sc_hd__a211o_1 _08586_ (.A1(_03148_),
    .A2(_03199_),
    .B1(_03206_),
    .C1(_02868_),
    .X(_03207_));
 sky130_fd_sc_hd__nand2_1 _08587_ (.A(_03166_),
    .B(_03207_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3_2 _08588_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03133_),
    .C(_03152_),
    .X(_03208_));
 sky130_fd_sc_hd__nor2_1 _08589_ (.A(_01971_),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__a221o_1 _08590_ (.A1(_01762_),
    .A2(_03208_),
    .B1(_03209_),
    .B2(net3236),
    .C1(_00209_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _08591_ (.A1(_01771_),
    .A2(_03208_),
    .B1(_03209_),
    .B2(net3143),
    .C1(_02872_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _08592_ (.A1(_01850_),
    .A2(_03208_),
    .B1(_03209_),
    .B2(net3260),
    .C1(_01973_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__mux4_1 _08593_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(_00792_),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A3(_00793_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .S1(net4154),
    .X(_03210_));
 sky130_fd_sc_hd__inv_2 _08594_ (.A(net3714),
    .Y(_03211_));
 sky130_fd_sc_hd__mux4_1 _08595_ (.A0(_00788_),
    .A1(_01060_),
    .A2(_01143_),
    .A3(_01059_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .S1(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__inv_2 _08596_ (.A(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__inv_2 _08597_ (.A(net3684),
    .Y(_03214_));
 sky130_fd_sc_hd__mux2_1 _08598_ (.A0(_03210_),
    .A1(_03213_),
    .S(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__clkbuf_1 _08599_ (.A(_03215_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ));
 sky130_fd_sc_hd__mux4_1 _08600_ (.A0(_01056_),
    .A1(_01059_),
    .A2(_00788_),
    .A3(_01061_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .X(_03216_));
 sky130_fd_sc_hd__clkinv_2 _08601_ (.A(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__mux4_1 _08602_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A3(_00793_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .X(_03218_));
 sky130_fd_sc_hd__mux2_1 _08603_ (.A0(_03217_),
    .A1(_03218_),
    .S(net3691),
    .X(_03219_));
 sky130_fd_sc_hd__clkbuf_1 _08604_ (.A(_03219_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ));
 sky130_fd_sc_hd__mux4_1 _08605_ (.A0(_00784_),
    .A1(_00786_),
    .A2(_00788_),
    .A3(_00789_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .X(_03220_));
 sky130_fd_sc_hd__clkinv_2 _08606_ (.A(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__mux4_1 _08607_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(_00792_),
    .A3(_00793_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(_03222_));
 sky130_fd_sc_hd__mux2_1 _08608_ (.A0(_03221_),
    .A1(_03222_),
    .S(net3707),
    .X(_03223_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08609_ (.A(_03223_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ));
 sky130_fd_sc_hd__mux4_1 _08610_ (.A0(_01227_),
    .A1(_01229_),
    .A2(_01059_),
    .A3(_01061_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .X(_03224_));
 sky130_fd_sc_hd__clkinv_2 _08611_ (.A(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__mux4_1 _08612_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A2(_00792_),
    .A3(_00793_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_1 _08613_ (.A0(_03225_),
    .A1(_03226_),
    .S(net3403),
    .X(_03227_));
 sky130_fd_sc_hd__clkbuf_1 _08614_ (.A(_03227_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ));
 sky130_fd_sc_hd__nor2_1 _08615_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ),
    .B(_02310_),
    .Y(_03228_));
 sky130_fd_sc_hd__mux2_1 _08616_ (.A0(_03104_),
    .A1(_03228_),
    .S(_01863_),
    .X(_03229_));
 sky130_fd_sc_hd__clkbuf_1 _08617_ (.A(_03229_),
    .X(_00005_));
 sky130_fd_sc_hd__nand3b_2 _08618_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .C(_01878_),
    .Y(_03230_));
 sky130_fd_sc_hd__or3_1 _08619_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_03231_));
 sky130_fd_sc_hd__or2_1 _08620_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_03231_),
    .X(_03232_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08621_ (.A(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__o21a_1 _08622_ (.A1(_03230_),
    .A2(_03233_),
    .B1(_03013_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_1 _08623_ (.A0(_03109_),
    .A1(net3325),
    .S(_03234_),
    .X(_03235_));
 sky130_fd_sc_hd__clkbuf_1 _08624_ (.A(_03235_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _08625_ (.A0(_03116_),
    .A1(net3358),
    .S(_03234_),
    .X(_03236_));
 sky130_fd_sc_hd__clkbuf_1 _08626_ (.A(_03236_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _08627_ (.A0(_03118_),
    .A1(net3299),
    .S(_03234_),
    .X(_03237_));
 sky130_fd_sc_hd__clkbuf_1 _08628_ (.A(_03237_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _08629_ (.A0(_03018_),
    .A1(net3480),
    .S(_03234_),
    .X(_03238_));
 sky130_fd_sc_hd__clkbuf_1 _08630_ (.A(_03238_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__clkbuf_2 _08631_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .X(_03239_));
 sky130_fd_sc_hd__inv_2 _08632_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .Y(_03240_));
 sky130_fd_sc_hd__or4_1 _08633_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_03239_),
    .C(_03240_),
    .D(_03230_),
    .X(_03241_));
 sky130_fd_sc_hd__o21a_2 _08634_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .A2(_03241_),
    .B1(_03013_),
    .X(_03242_));
 sky130_fd_sc_hd__mux2_1 _08635_ (.A0(_03109_),
    .A1(net3562),
    .S(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__clkbuf_1 _08636_ (.A(_03243_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _08637_ (.A0(_03116_),
    .A1(net3343),
    .S(_03242_),
    .X(_03244_));
 sky130_fd_sc_hd__clkbuf_1 _08638_ (.A(_03244_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _08639_ (.A0(_03118_),
    .A1(net3755),
    .S(_03242_),
    .X(_03245_));
 sky130_fd_sc_hd__clkbuf_1 _08640_ (.A(_03245_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__buf_4 _08641_ (.A(_00191_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _08642_ (.A0(_03246_),
    .A1(net3751),
    .S(_03242_),
    .X(_03247_));
 sky130_fd_sc_hd__clkbuf_1 _08643_ (.A(_03247_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _08644_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .Y(_03248_));
 sky130_fd_sc_hd__or3_2 _08645_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(_03248_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_03249_));
 sky130_fd_sc_hd__and3b_1 _08646_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .C(_00311_),
    .X(_03250_));
 sky130_fd_sc_hd__nand2_1 _08647_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_03231_),
    .Y(_03251_));
 sky130_fd_sc_hd__and2_1 _08648_ (.A(_03233_),
    .B(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__nand2_1 _08649_ (.A(_03250_),
    .B(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__nand2_1 _08650_ (.A(_00170_),
    .B(_03233_),
    .Y(_03254_));
 sky130_fd_sc_hd__or3_1 _08651_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_03230_),
    .C(_03249_),
    .X(_03255_));
 sky130_fd_sc_hd__nand2_1 _08652_ (.A(net3560),
    .B(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__o31a_1 _08653_ (.A1(_03249_),
    .A2(_03253_),
    .A3(_03254_),
    .B1(_03256_),
    .X(_03257_));
 sky130_fd_sc_hd__o21ai_1 _08654_ (.A1(_03141_),
    .A2(_03257_),
    .B1(_02978_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_1 _08655_ (.A(_00211_),
    .B(_03233_),
    .Y(_03258_));
 sky130_fd_sc_hd__nand2_1 _08656_ (.A(net3496),
    .B(_03255_),
    .Y(_03259_));
 sky130_fd_sc_hd__o31a_1 _08657_ (.A1(_03249_),
    .A2(_03253_),
    .A3(_03258_),
    .B1(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__o21ai_1 _08658_ (.A1(_03141_),
    .A2(_03260_),
    .B1(_02714_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__nand2_1 _08659_ (.A(_02573_),
    .B(_03233_),
    .Y(_03261_));
 sky130_fd_sc_hd__nand2_1 _08660_ (.A(net3718),
    .B(_03255_),
    .Y(_03262_));
 sky130_fd_sc_hd__o31a_1 _08661_ (.A1(_03249_),
    .A2(_03253_),
    .A3(_03261_),
    .B1(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__o21ai_1 _08662_ (.A1(_03141_),
    .A2(_03263_),
    .B1(_02740_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__clkbuf_4 _08663_ (.A(_01764_),
    .X(_03264_));
 sky130_fd_sc_hd__nand2_1 _08664_ (.A(_01452_),
    .B(_03233_),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2_1 _08665_ (.A(net3754),
    .B(_03255_),
    .Y(_03266_));
 sky130_fd_sc_hd__o31a_1 _08666_ (.A1(_03249_),
    .A2(_03253_),
    .A3(_03265_),
    .B1(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__o21ai_1 _08667_ (.A1(_03264_),
    .A2(_03267_),
    .B1(_02928_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_1 _08668_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_03230_),
    .Y(_03268_));
 sky130_fd_sc_hd__and3b_1 _08669_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_03269_));
 sky130_fd_sc_hd__a21oi_2 _08670_ (.A1(_03268_),
    .A2(_03269_),
    .B1(_02686_),
    .Y(_03270_));
 sky130_fd_sc_hd__mux2_1 _08671_ (.A0(_03109_),
    .A1(net3456),
    .S(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__clkbuf_1 _08672_ (.A(_03271_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _08673_ (.A0(_03116_),
    .A1(net3396),
    .S(_03270_),
    .X(_03272_));
 sky130_fd_sc_hd__clkbuf_1 _08674_ (.A(_03272_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _08675_ (.A0(_03118_),
    .A1(net3448),
    .S(_03270_),
    .X(_03273_));
 sky130_fd_sc_hd__clkbuf_1 _08676_ (.A(_03273_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _08677_ (.A0(_03246_),
    .A1(net3357),
    .S(_03270_),
    .X(_03274_));
 sky130_fd_sc_hd__clkbuf_1 _08678_ (.A(_03274_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4_1 _08679_ (.A(_03239_),
    .B(_03248_),
    .C(_03240_),
    .D(_03268_),
    .X(_03275_));
 sky130_fd_sc_hd__clkbuf_2 _08680_ (.A(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__nand2_1 _08681_ (.A(_03254_),
    .B(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__or2_1 _08682_ (.A(net4129),
    .B(_03276_),
    .X(_03278_));
 sky130_fd_sc_hd__a31o_1 _08683_ (.A1(_03085_),
    .A2(_03277_),
    .A3(_03278_),
    .B1(_02711_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _08684_ (.A(_03258_),
    .B(_03276_),
    .Y(_03279_));
 sky130_fd_sc_hd__or2_1 _08685_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .B(_03276_),
    .X(_03280_));
 sky130_fd_sc_hd__a31o_1 _08686_ (.A1(_03085_),
    .A2(_03279_),
    .A3(_03280_),
    .B1(_03050_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__clkbuf_4 _08687_ (.A(_00195_),
    .X(_03281_));
 sky130_fd_sc_hd__nand2_1 _08688_ (.A(_03261_),
    .B(_03276_),
    .Y(_03282_));
 sky130_fd_sc_hd__or2_1 _08689_ (.A(net4208),
    .B(_03276_),
    .X(_03283_));
 sky130_fd_sc_hd__a31o_1 _08690_ (.A1(_03281_),
    .A2(_03282_),
    .A3(_03283_),
    .B1(_01851_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _08691_ (.A(net4019),
    .B(_03276_),
    .Y(_03284_));
 sky130_fd_sc_hd__a211o_1 _08692_ (.A1(_03265_),
    .A2(_03276_),
    .B1(_03284_),
    .C1(_02868_),
    .X(_03285_));
 sky130_fd_sc_hd__nand2_1 _08693_ (.A(_03166_),
    .B(_03285_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _08694_ (.A1(_03239_),
    .A2(_03248_),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .A4(_03268_),
    .B1(_02946_),
    .X(_03286_));
 sky130_fd_sc_hd__mux2_1 _08695_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .A1(_03169_),
    .S(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__clkbuf_1 _08696_ (.A(_03287_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _08697_ (.A0(net4171),
    .A1(_03172_),
    .S(_03286_),
    .X(_03288_));
 sky130_fd_sc_hd__clkbuf_1 _08698_ (.A(_03288_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _08699_ (.A0(net3836),
    .A1(_03174_),
    .S(_03286_),
    .X(_03289_));
 sky130_fd_sc_hd__clkbuf_1 _08700_ (.A(_03289_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _08701_ (.A0(net3205),
    .A1(_02951_),
    .S(_03286_),
    .X(_03290_));
 sky130_fd_sc_hd__clkbuf_1 _08702_ (.A(_03290_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_1 _08703_ (.A(_03239_),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .C(_03240_),
    .D(_03268_),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _08704_ (.A0(_02384_),
    .A1(_03254_),
    .S(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__o21ai_1 _08705_ (.A1(_03264_),
    .A2(_03292_),
    .B1(_02978_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _08706_ (.A0(_02385_),
    .A1(_03258_),
    .S(_03291_),
    .X(_03293_));
 sky130_fd_sc_hd__o21ai_1 _08707_ (.A1(_03264_),
    .A2(_03293_),
    .B1(_02714_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _08708_ (.A0(_02389_),
    .A1(_03261_),
    .S(_03291_),
    .X(_03294_));
 sky130_fd_sc_hd__o21ai_1 _08709_ (.A1(_03264_),
    .A2(_03294_),
    .B1(_02740_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _08710_ (.A0(_02380_),
    .A1(_03265_),
    .S(_03291_),
    .X(_03295_));
 sky130_fd_sc_hd__o21ai_1 _08711_ (.A1(_03264_),
    .A2(_03295_),
    .B1(_02928_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _08712_ (.A1(_03239_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .A4(_03268_),
    .B1(_02946_),
    .X(_03296_));
 sky130_fd_sc_hd__mux2_1 _08713_ (.A0(net3610),
    .A1(_03169_),
    .S(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__clkbuf_1 _08714_ (.A(_03297_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _08715_ (.A0(net4186),
    .A1(_03172_),
    .S(_03296_),
    .X(_03298_));
 sky130_fd_sc_hd__clkbuf_1 _08716_ (.A(_03298_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _08717_ (.A0(net3935),
    .A1(_03174_),
    .S(_03296_),
    .X(_03299_));
 sky130_fd_sc_hd__clkbuf_1 _08718_ (.A(_03299_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _08719_ (.A0(net3889),
    .A1(_02951_),
    .S(_03296_),
    .X(_03300_));
 sky130_fd_sc_hd__clkbuf_1 _08720_ (.A(_03300_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _08721_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .Y(_03301_));
 sky130_fd_sc_hd__o31a_1 _08722_ (.A1(_03301_),
    .A2(_03230_),
    .A3(_03231_),
    .B1(_02847_),
    .X(_03302_));
 sky130_fd_sc_hd__mux2_1 _08723_ (.A0(_03109_),
    .A1(net3775),
    .S(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__clkbuf_1 _08724_ (.A(_03303_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _08725_ (.A0(_03116_),
    .A1(net3442),
    .S(_03302_),
    .X(_03304_));
 sky130_fd_sc_hd__clkbuf_1 _08726_ (.A(_03304_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _08727_ (.A0(_03118_),
    .A1(net3698),
    .S(_03302_),
    .X(_03305_));
 sky130_fd_sc_hd__clkbuf_1 _08728_ (.A(_03305_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _08729_ (.A0(_03246_),
    .A1(net3981),
    .S(_03302_),
    .X(_03306_));
 sky130_fd_sc_hd__clkbuf_1 _08730_ (.A(_03306_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _08731_ (.A(_03230_),
    .B(_03252_),
    .X(_03307_));
 sky130_fd_sc_hd__o41a_2 _08732_ (.A1(_03239_),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .A3(_03240_),
    .A4(_03307_),
    .B1(_00407_),
    .X(_03308_));
 sky130_fd_sc_hd__mux2_1 _08733_ (.A0(_03109_),
    .A1(net3617),
    .S(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__clkbuf_1 _08734_ (.A(_03309_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _08735_ (.A0(_03116_),
    .A1(net3380),
    .S(_03308_),
    .X(_03310_));
 sky130_fd_sc_hd__clkbuf_1 _08736_ (.A(_03310_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _08737_ (.A0(_03118_),
    .A1(net3952),
    .S(_03308_),
    .X(_03311_));
 sky130_fd_sc_hd__clkbuf_1 _08738_ (.A(_03311_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _08739_ (.A0(_03246_),
    .A1(net3605),
    .S(_03308_),
    .X(_03312_));
 sky130_fd_sc_hd__clkbuf_1 _08740_ (.A(_03312_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _08741_ (.A(_03249_),
    .B(_03307_),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_1 _08742_ (.A(_03254_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__or2_1 _08743_ (.A(net4039),
    .B(_03313_),
    .X(_03315_));
 sky130_fd_sc_hd__buf_6 _08744_ (.A(_00208_),
    .X(_03316_));
 sky130_fd_sc_hd__a31o_1 _08745_ (.A1(_03281_),
    .A2(_03314_),
    .A3(_03315_),
    .B1(_03316_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__or2_1 _08746_ (.A(net3936),
    .B(_03313_),
    .X(_03317_));
 sky130_fd_sc_hd__nand2_1 _08747_ (.A(_03258_),
    .B(_03313_),
    .Y(_03318_));
 sky130_fd_sc_hd__a31o_1 _08748_ (.A1(_03281_),
    .A2(_03317_),
    .A3(_03318_),
    .B1(_03050_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__or2_1 _08749_ (.A(net3523),
    .B(_03313_),
    .X(_03319_));
 sky130_fd_sc_hd__nand2_1 _08750_ (.A(_03261_),
    .B(_03313_),
    .Y(_03320_));
 sky130_fd_sc_hd__a31o_1 _08751_ (.A1(_03281_),
    .A2(_03319_),
    .A3(_03320_),
    .B1(_01851_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__mux2_1 _08752_ (.A0(_02830_),
    .A1(_03265_),
    .S(_03313_),
    .X(_03321_));
 sky130_fd_sc_hd__clkbuf_8 _08753_ (.A(_00226_),
    .X(_03322_));
 sky130_fd_sc_hd__o21ai_1 _08754_ (.A1(_03264_),
    .A2(_03321_),
    .B1(_03322_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3_2 _08755_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_03250_),
    .C(_03269_),
    .X(_03323_));
 sky130_fd_sc_hd__nor2_1 _08756_ (.A(_01971_),
    .B(_03323_),
    .Y(_03324_));
 sky130_fd_sc_hd__a221o_1 _08757_ (.A1(_00288_),
    .A2(_03323_),
    .B1(_03324_),
    .B2(net3382),
    .C1(_00209_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _08758_ (.A1(_00293_),
    .A2(_03323_),
    .B1(_03324_),
    .B2(net3173),
    .C1(_02872_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _08759_ (.A1(_00295_),
    .A2(_03323_),
    .B1(_03324_),
    .B2(net3138),
    .C1(_01973_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__mux4_1 _08760_ (.A0(_01143_),
    .A1(_01058_),
    .A2(_00788_),
    .A3(_01061_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .X(_03325_));
 sky130_fd_sc_hd__clkinv_2 _08761_ (.A(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__mux4_1 _08762_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A3(_00793_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .X(_03327_));
 sky130_fd_sc_hd__mux2_1 _08763_ (.A0(_03326_),
    .A1(_03327_),
    .S(net3337),
    .X(_03328_));
 sky130_fd_sc_hd__clkbuf_1 _08764_ (.A(net3338),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ));
 sky130_fd_sc_hd__mux4_1 _08765_ (.A0(_01056_),
    .A1(_01058_),
    .A2(_00788_),
    .A3(_01061_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .X(_03329_));
 sky130_fd_sc_hd__clkinv_2 _08766_ (.A(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__mux4_1 _08767_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .X(_03331_));
 sky130_fd_sc_hd__mux2_1 _08768_ (.A0(_03330_),
    .A1(_03331_),
    .S(net3477),
    .X(_03332_));
 sky130_fd_sc_hd__clkbuf_1 _08769_ (.A(_03332_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ));
 sky130_fd_sc_hd__mux4_1 _08770_ (.A0(_00784_),
    .A1(_00786_),
    .A2(_00787_),
    .A3(_00789_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .X(_03333_));
 sky130_fd_sc_hd__clkinv_2 _08771_ (.A(_03333_),
    .Y(_03334_));
 sky130_fd_sc_hd__mux4_1 _08772_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(_00792_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _08773_ (.A0(_03334_),
    .A1(_03335_),
    .S(net3468),
    .X(_03336_));
 sky130_fd_sc_hd__clkbuf_1 _08774_ (.A(_03336_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ));
 sky130_fd_sc_hd__mux4_1 _08775_ (.A0(_01227_),
    .A1(_01229_),
    .A2(_01059_),
    .A3(_01061_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .X(_03337_));
 sky130_fd_sc_hd__clkinv_2 _08776_ (.A(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__mux4_1 _08777_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A2(_00792_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_1 _08778_ (.A0(_03338_),
    .A1(_03339_),
    .S(net3630),
    .X(_03340_));
 sky130_fd_sc_hd__clkbuf_1 _08779_ (.A(_03340_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ));
 sky130_fd_sc_hd__a22o_1 _08780_ (.A1(_02394_),
    .A2(_02398_),
    .B1(_02400_),
    .B2(_02404_),
    .X(_03341_));
 sky130_fd_sc_hd__and2_1 _08781_ (.A(_01858_),
    .B(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_1 _08782_ (.A0(_03228_),
    .A1(_03342_),
    .S(_01863_),
    .X(_03343_));
 sky130_fd_sc_hd__clkbuf_1 _08783_ (.A(_03343_),
    .X(_00006_));
 sky130_fd_sc_hd__buf_4 _08784_ (.A(_00171_),
    .X(_03344_));
 sky130_fd_sc_hd__nand3b_2 _08785_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .C(_01878_),
    .Y(_03345_));
 sky130_fd_sc_hd__or3_1 _08786_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_03346_));
 sky130_fd_sc_hd__or2_1 _08787_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_03346_),
    .X(_03347_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08788_ (.A(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__o21a_2 _08789_ (.A1(_03345_),
    .A2(_03348_),
    .B1(_03013_),
    .X(_03349_));
 sky130_fd_sc_hd__mux2_1 _08790_ (.A0(_03344_),
    .A1(net3414),
    .S(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__clkbuf_1 _08791_ (.A(_03350_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__buf_4 _08792_ (.A(_00184_),
    .X(_03351_));
 sky130_fd_sc_hd__mux2_1 _08793_ (.A0(_03351_),
    .A1(net3413),
    .S(_03349_),
    .X(_03352_));
 sky130_fd_sc_hd__clkbuf_1 _08794_ (.A(_03352_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__buf_4 _08795_ (.A(_00551_),
    .X(_03353_));
 sky130_fd_sc_hd__mux2_1 _08796_ (.A0(_03353_),
    .A1(net3580),
    .S(_03349_),
    .X(_03354_));
 sky130_fd_sc_hd__clkbuf_1 _08797_ (.A(_03354_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _08798_ (.A0(_03246_),
    .A1(net3673),
    .S(_03349_),
    .X(_03355_));
 sky130_fd_sc_hd__clkbuf_1 _08799_ (.A(_03355_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _08800_ (.A(net4168),
    .X(_03356_));
 sky130_fd_sc_hd__clkbuf_2 _08801_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .X(_03357_));
 sky130_fd_sc_hd__inv_2 _08802_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .Y(_03358_));
 sky130_fd_sc_hd__or4_1 _08803_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_03357_),
    .C(_03358_),
    .D(_03345_),
    .X(_03359_));
 sky130_fd_sc_hd__o21a_2 _08804_ (.A1(_03356_),
    .A2(_03359_),
    .B1(_03013_),
    .X(_03360_));
 sky130_fd_sc_hd__mux2_1 _08805_ (.A0(_03344_),
    .A1(net3316),
    .S(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__clkbuf_1 _08806_ (.A(_03361_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _08807_ (.A0(_03351_),
    .A1(net3586),
    .S(_03360_),
    .X(_03362_));
 sky130_fd_sc_hd__clkbuf_1 _08808_ (.A(_03362_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _08809_ (.A0(_03353_),
    .A1(net3578),
    .S(_03360_),
    .X(_03363_));
 sky130_fd_sc_hd__clkbuf_1 _08810_ (.A(_03363_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _08811_ (.A0(_03246_),
    .A1(net3339),
    .S(_03360_),
    .X(_03364_));
 sky130_fd_sc_hd__clkbuf_1 _08812_ (.A(_03364_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _08813_ (.A(_03356_),
    .Y(_03365_));
 sky130_fd_sc_hd__or3_2 _08814_ (.A(_03357_),
    .B(_03365_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_03366_));
 sky130_fd_sc_hd__and3b_1 _08815_ (.A_N(\c.genblk1.genblk1.subs.cs[1].c.cfgd ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .C(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_2 _08816_ (.A(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__nand2_1 _08817_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_03346_),
    .Y(_03369_));
 sky130_fd_sc_hd__and2_1 _08818_ (.A(_03348_),
    .B(_03369_),
    .X(_03370_));
 sky130_fd_sc_hd__nand2_1 _08819_ (.A(_03368_),
    .B(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand2_1 _08820_ (.A(_00170_),
    .B(_03348_),
    .Y(_03372_));
 sky130_fd_sc_hd__or3_1 _08821_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_03345_),
    .C(_03366_),
    .X(_03373_));
 sky130_fd_sc_hd__nand2_1 _08822_ (.A(net3850),
    .B(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__o31a_1 _08823_ (.A1(_03366_),
    .A2(_03371_),
    .A3(_03372_),
    .B1(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__o21ai_1 _08824_ (.A1(_03264_),
    .A2(_03375_),
    .B1(_02978_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_1 _08825_ (.A(_00211_),
    .B(_03348_),
    .Y(_03376_));
 sky130_fd_sc_hd__nand2_1 _08826_ (.A(net3485),
    .B(_03373_),
    .Y(_03377_));
 sky130_fd_sc_hd__o31a_1 _08827_ (.A1(_03366_),
    .A2(_03371_),
    .A3(_03376_),
    .B1(_03377_),
    .X(_03378_));
 sky130_fd_sc_hd__buf_4 _08828_ (.A(_00305_),
    .X(_03379_));
 sky130_fd_sc_hd__o21ai_1 _08829_ (.A1(_03264_),
    .A2(_03378_),
    .B1(_03379_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__nand2_1 _08830_ (.A(_02573_),
    .B(_03348_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand2_1 _08831_ (.A(net3747),
    .B(_03373_),
    .Y(_03381_));
 sky130_fd_sc_hd__o31a_1 _08832_ (.A1(_03366_),
    .A2(_03371_),
    .A3(_03380_),
    .B1(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__o21ai_1 _08833_ (.A1(_03264_),
    .A2(_03382_),
    .B1(_00251_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__nand2_1 _08834_ (.A(_00264_),
    .B(_03348_),
    .Y(_03383_));
 sky130_fd_sc_hd__nand2_1 _08835_ (.A(net3393),
    .B(_03373_),
    .Y(_03384_));
 sky130_fd_sc_hd__o31a_1 _08836_ (.A1(_03366_),
    .A2(_03371_),
    .A3(_03383_),
    .B1(_03384_),
    .X(_03385_));
 sky130_fd_sc_hd__o21ai_1 _08837_ (.A1(_03264_),
    .A2(_03385_),
    .B1(_03322_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _08838_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_03345_),
    .Y(_03386_));
 sky130_fd_sc_hd__and3b_1 _08839_ (.A_N(_03357_),
    .B(_03356_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_03387_));
 sky130_fd_sc_hd__a21oi_4 _08840_ (.A1(_03386_),
    .A2(_03387_),
    .B1(_02686_),
    .Y(_03388_));
 sky130_fd_sc_hd__mux2_1 _08841_ (.A0(_03344_),
    .A1(net3546),
    .S(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_1 _08842_ (.A(_03389_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _08843_ (.A0(_03351_),
    .A1(net3582),
    .S(_03388_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_1 _08844_ (.A(_03390_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _08845_ (.A0(_03353_),
    .A1(net3320),
    .S(_03388_),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_1 _08846_ (.A(_03391_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _08847_ (.A0(_03246_),
    .A1(net3441),
    .S(_03388_),
    .X(_03392_));
 sky130_fd_sc_hd__clkbuf_1 _08848_ (.A(_03392_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4_1 _08849_ (.A(_03357_),
    .B(_03365_),
    .C(_03358_),
    .D(_03386_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_2 _08850_ (.A(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__nand2_1 _08851_ (.A(_03372_),
    .B(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__or2_1 _08852_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .B(_03394_),
    .X(_03396_));
 sky130_fd_sc_hd__a31o_1 _08853_ (.A1(_03281_),
    .A2(_03395_),
    .A3(_03396_),
    .B1(_03316_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _08854_ (.A(_03376_),
    .B(_03394_),
    .Y(_03397_));
 sky130_fd_sc_hd__or2_1 _08855_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .B(_03394_),
    .X(_03398_));
 sky130_fd_sc_hd__a31o_1 _08856_ (.A1(_03281_),
    .A2(_03397_),
    .A3(_03398_),
    .B1(_03050_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _08857_ (.A(_03380_),
    .B(_03394_),
    .Y(_03399_));
 sky130_fd_sc_hd__or2_1 _08858_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .B(_03394_),
    .X(_03400_));
 sky130_fd_sc_hd__a31o_1 _08859_ (.A1(_03281_),
    .A2(_03399_),
    .A3(_03400_),
    .B1(_01851_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _08860_ (.A(net4183),
    .B(_03394_),
    .Y(_03401_));
 sky130_fd_sc_hd__a211o_1 _08861_ (.A1(_03383_),
    .A2(_03394_),
    .B1(_03401_),
    .C1(_02868_),
    .X(_03402_));
 sky130_fd_sc_hd__nand2_1 _08862_ (.A(_03166_),
    .B(_03402_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _08863_ (.A1(_03357_),
    .A2(_03365_),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .A4(_03386_),
    .B1(_02946_),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_1 _08864_ (.A0(net4009),
    .A1(_03169_),
    .S(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_1 _08865_ (.A(_03404_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _08866_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .A1(_03172_),
    .S(_03403_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_1 _08867_ (.A(_03405_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _08868_ (.A0(net4003),
    .A1(_03174_),
    .S(_03403_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_1 _08869_ (.A(_03406_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _08870_ (.A0(net3932),
    .A1(_02951_),
    .S(_03403_),
    .X(_03407_));
 sky130_fd_sc_hd__clkbuf_1 _08871_ (.A(_03407_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__buf_4 _08872_ (.A(_01764_),
    .X(_03408_));
 sky130_fd_sc_hd__and4_1 _08873_ (.A(_03357_),
    .B(_03356_),
    .C(_03358_),
    .D(_03386_),
    .X(_03409_));
 sky130_fd_sc_hd__mux2_1 _08874_ (.A0(_02425_),
    .A1(_03372_),
    .S(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__o21ai_1 _08875_ (.A1(_03408_),
    .A2(_03410_),
    .B1(_02978_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _08876_ (.A0(_02426_),
    .A1(_03376_),
    .S(_03409_),
    .X(_03411_));
 sky130_fd_sc_hd__o21ai_1 _08877_ (.A1(_03408_),
    .A2(_03411_),
    .B1(_03379_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _08878_ (.A0(_02430_),
    .A1(_03380_),
    .S(_03409_),
    .X(_03412_));
 sky130_fd_sc_hd__o21ai_1 _08879_ (.A1(_03408_),
    .A2(_03412_),
    .B1(_00251_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _08880_ (.A0(_02420_),
    .A1(_03383_),
    .S(_03409_),
    .X(_03413_));
 sky130_fd_sc_hd__o21ai_1 _08881_ (.A1(_03408_),
    .A2(_03413_),
    .B1(_03322_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _08882_ (.A1(_03357_),
    .A2(_03356_),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .A4(_03386_),
    .B1(_02946_),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_1 _08883_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .A1(_03169_),
    .S(_03414_),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_1 _08884_ (.A(_03415_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _08885_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A1(_03172_),
    .S(_03414_),
    .X(_03416_));
 sky130_fd_sc_hd__clkbuf_1 _08886_ (.A(_03416_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _08887_ (.A0(net3778),
    .A1(_03174_),
    .S(_03414_),
    .X(_03417_));
 sky130_fd_sc_hd__clkbuf_1 _08888_ (.A(_03417_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _08889_ (.A0(net4135),
    .A1(_02951_),
    .S(_03414_),
    .X(_03418_));
 sky130_fd_sc_hd__clkbuf_1 _08890_ (.A(_03418_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _08891_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .Y(_03419_));
 sky130_fd_sc_hd__o31a_2 _08892_ (.A1(_03419_),
    .A2(_03345_),
    .A3(_03346_),
    .B1(_02847_),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_1 _08893_ (.A0(_03344_),
    .A1(net3131),
    .S(_03420_),
    .X(_03421_));
 sky130_fd_sc_hd__clkbuf_1 _08894_ (.A(net3132),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _08895_ (.A0(_03351_),
    .A1(net3705),
    .S(_03420_),
    .X(_03422_));
 sky130_fd_sc_hd__clkbuf_1 _08896_ (.A(_03422_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _08897_ (.A0(_03353_),
    .A1(net3942),
    .S(_03420_),
    .X(_03423_));
 sky130_fd_sc_hd__clkbuf_1 _08898_ (.A(_03423_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _08899_ (.A0(_03246_),
    .A1(net3313),
    .S(_03420_),
    .X(_03424_));
 sky130_fd_sc_hd__clkbuf_1 _08900_ (.A(_03424_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _08901_ (.A(_03345_),
    .B(_03370_),
    .X(_03425_));
 sky130_fd_sc_hd__o41a_2 _08902_ (.A1(_03357_),
    .A2(_03356_),
    .A3(_03358_),
    .A4(_03425_),
    .B1(_00407_),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_1 _08903_ (.A0(_03344_),
    .A1(net3838),
    .S(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__clkbuf_1 _08904_ (.A(_03427_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _08905_ (.A0(_03351_),
    .A1(net3720),
    .S(_03426_),
    .X(_03428_));
 sky130_fd_sc_hd__clkbuf_1 _08906_ (.A(_03428_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _08907_ (.A0(_03353_),
    .A1(net3839),
    .S(_03426_),
    .X(_03429_));
 sky130_fd_sc_hd__clkbuf_1 _08908_ (.A(_03429_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _08909_ (.A0(_03246_),
    .A1(net3541),
    .S(_03426_),
    .X(_03430_));
 sky130_fd_sc_hd__clkbuf_1 _08910_ (.A(_03430_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _08911_ (.A(_03366_),
    .B(_03425_),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_1 _08912_ (.A(_03372_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__or2_1 _08913_ (.A(net3780),
    .B(_03431_),
    .X(_03433_));
 sky130_fd_sc_hd__a31o_1 _08914_ (.A1(_03281_),
    .A2(_03432_),
    .A3(_03433_),
    .B1(_03316_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__or2_1 _08915_ (.A(net4059),
    .B(_03431_),
    .X(_03434_));
 sky130_fd_sc_hd__nand2_1 _08916_ (.A(_03376_),
    .B(_03431_),
    .Y(_03435_));
 sky130_fd_sc_hd__a31o_1 _08917_ (.A1(_03281_),
    .A2(_03434_),
    .A3(_03435_),
    .B1(_03050_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__nand2_1 _08918_ (.A(_03380_),
    .B(_03431_),
    .Y(_03436_));
 sky130_fd_sc_hd__or2_1 _08919_ (.A(net3160),
    .B(_03431_),
    .X(_03437_));
 sky130_fd_sc_hd__a31o_1 _08920_ (.A1(_03281_),
    .A2(_03436_),
    .A3(_03437_),
    .B1(_01851_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__nor2_1 _08921_ (.A(net3979),
    .B(_03431_),
    .Y(_03438_));
 sky130_fd_sc_hd__a211o_1 _08922_ (.A1(_03383_),
    .A2(_03431_),
    .B1(_03438_),
    .C1(_02868_),
    .X(_03439_));
 sky130_fd_sc_hd__nand2_1 _08923_ (.A(_03166_),
    .B(_03439_),
    .Y(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3_2 _08924_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_03368_),
    .C(_03387_),
    .X(_03440_));
 sky130_fd_sc_hd__nor2_1 _08925_ (.A(_01971_),
    .B(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__a221o_1 _08926_ (.A1(_00288_),
    .A2(_03440_),
    .B1(_03441_),
    .B2(net3657),
    .C1(_00209_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _08927_ (.A1(_00293_),
    .A2(_03440_),
    .B1(_03441_),
    .B2(net3167),
    .C1(_02872_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _08928_ (.A1(_00295_),
    .A2(_03440_),
    .B1(_03441_),
    .B2(net3212),
    .C1(_00221_),
    .X(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__inv_2 _08929_ (.A(net3695),
    .Y(_03442_));
 sky130_fd_sc_hd__mux4_1 _08930_ (.A0(_00788_),
    .A1(_01060_),
    .A2(_01143_),
    .A3(_01059_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ),
    .S1(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__clkinv_2 _08931_ (.A(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__mux4_1 _08932_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ),
    .S1(net4218),
    .X(_03445_));
 sky130_fd_sc_hd__mux2_1 _08933_ (.A0(_03444_),
    .A1(_03445_),
    .S(net3312),
    .X(_03446_));
 sky130_fd_sc_hd__clkbuf_1 _08934_ (.A(_03446_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ));
 sky130_fd_sc_hd__inv_2 _08935_ (.A(net3694),
    .Y(_03447_));
 sky130_fd_sc_hd__mux4_1 _08936_ (.A0(_01059_),
    .A1(_01056_),
    .A2(_01061_),
    .A3(_00788_),
    .S0(_03447_),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .X(_03448_));
 sky130_fd_sc_hd__clkinv_2 _08937_ (.A(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__mux4_1 _08938_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .X(_03450_));
 sky130_fd_sc_hd__mux2_1 _08939_ (.A0(_03449_),
    .A1(_03450_),
    .S(net3589),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_1 _08940_ (.A(_03451_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ));
 sky130_fd_sc_hd__mux4_1 _08941_ (.A0(_00784_),
    .A1(_00786_),
    .A2(_00787_),
    .A3(_00789_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .X(_03452_));
 sky130_fd_sc_hd__clkinv_2 _08942_ (.A(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__mux4_1 _08943_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ),
    .A2(_00792_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ),
    .X(_03454_));
 sky130_fd_sc_hd__mux2_1 _08944_ (.A0(_03453_),
    .A1(_03454_),
    .S(net3438),
    .X(_03455_));
 sky130_fd_sc_hd__clkbuf_1 _08945_ (.A(_03455_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ));
 sky130_fd_sc_hd__mux4_1 _08946_ (.A0(_01227_),
    .A1(_01229_),
    .A2(_01059_),
    .A3(_01061_),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .X(_03456_));
 sky130_fd_sc_hd__clkinv_2 _08947_ (.A(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__mux4_1 _08948_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ),
    .A2(_00792_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ),
    .S0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .S1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .X(_03458_));
 sky130_fd_sc_hd__mux2_1 _08949_ (.A0(_03457_),
    .A1(_03458_),
    .S(net3412),
    .X(_03459_));
 sky130_fd_sc_hd__clkbuf_1 _08950_ (.A(_03459_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ));
 sky130_fd_sc_hd__mux2_1 _08951_ (.A0(_03103_),
    .A1(_03342_),
    .S(_02524_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_1 _08952_ (.A(_03460_),
    .X(_00007_));
 sky130_fd_sc_hd__clkbuf_4 _08953_ (.A(_01580_),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_4 _08954_ (.A(_01673_),
    .X(_03462_));
 sky130_fd_sc_hd__buf_4 _08955_ (.A(_01759_),
    .X(_03463_));
 sky130_fd_sc_hd__buf_4 _08956_ (.A(_01849_),
    .X(_03464_));
 sky130_fd_sc_hd__mux4_1 _08957_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[36] ),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_4 _08958_ (.A(net11),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_4 _08959_ (.A(net18),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_4 _08960_ (.A(net19),
    .X(_03468_));
 sky130_fd_sc_hd__clkbuf_4 _08961_ (.A(net20),
    .X(_03469_));
 sky130_fd_sc_hd__mux4_1 _08962_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[36] ),
    .X(_03470_));
 sky130_fd_sc_hd__nor2_1 _08963_ (.A(_00307_),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__a211o_1 _08964_ (.A1(_00307_),
    .A2(_03465_),
    .B1(_03471_),
    .C1(_00303_),
    .X(_03472_));
 sky130_fd_sc_hd__clkbuf_4 _08965_ (.A(_01311_),
    .X(_03473_));
 sky130_fd_sc_hd__clkbuf_4 _08966_ (.A(_01395_),
    .X(_03474_));
 sky130_fd_sc_hd__mux4_1 _08967_ (.A0(_00880_),
    .A1(_00972_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[36] ),
    .X(_03475_));
 sky130_fd_sc_hd__or3_1 _08968_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[37] ),
    .B(_00307_),
    .C(_03475_),
    .X(_03476_));
 sky130_fd_sc_hd__nor2_1 _08969_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[37] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[38] ),
    .Y(_03477_));
 sky130_fd_sc_hd__buf_2 _08970_ (.A(_02226_),
    .X(_03478_));
 sky130_fd_sc_hd__clkbuf_2 _08971_ (.A(_02320_),
    .X(_03479_));
 sky130_fd_sc_hd__clkbuf_2 _08972_ (.A(_02408_),
    .X(_03480_));
 sky130_fd_sc_hd__clkbuf_2 _08973_ (.A(_02491_),
    .X(_03481_));
 sky130_fd_sc_hd__mux4_1 _08974_ (.A0(_03478_),
    .A1(_03479_),
    .A2(_03480_),
    .A3(_03481_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[36] ),
    .X(_03482_));
 sky130_fd_sc_hd__a21oi_1 _08975_ (.A1(_03477_),
    .A2(_03482_),
    .B1(net3631),
    .Y(_03483_));
 sky130_fd_sc_hd__clkbuf_4 _08976_ (.A(net21),
    .X(_03484_));
 sky130_fd_sc_hd__clkbuf_4 _08977_ (.A(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__clkbuf_4 _08978_ (.A(net22),
    .X(_03486_));
 sky130_fd_sc_hd__clkbuf_4 _08979_ (.A(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__clkbuf_4 _08980_ (.A(net23),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_4 _08981_ (.A(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__clkbuf_4 _08982_ (.A(net24),
    .X(_03490_));
 sky130_fd_sc_hd__clkbuf_4 _08983_ (.A(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__mux4_1 _08984_ (.A0(_03485_),
    .A1(_03487_),
    .A2(_03489_),
    .A3(_03491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[36] ),
    .X(_03492_));
 sky130_fd_sc_hd__clkbuf_4 _08985_ (.A(net14),
    .X(_03493_));
 sky130_fd_sc_hd__clkbuf_4 _08986_ (.A(_03493_),
    .X(_03494_));
 sky130_fd_sc_hd__clkbuf_4 _08987_ (.A(net15),
    .X(_03495_));
 sky130_fd_sc_hd__clkbuf_4 _08988_ (.A(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__clkbuf_4 _08989_ (.A(net16),
    .X(_03497_));
 sky130_fd_sc_hd__clkbuf_4 _08990_ (.A(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__clkbuf_4 _08991_ (.A(net17),
    .X(_03499_));
 sky130_fd_sc_hd__clkbuf_4 _08992_ (.A(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__mux4_1 _08993_ (.A0(_03494_),
    .A1(_03496_),
    .A2(_03498_),
    .A3(_03500_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[36] ),
    .X(_03501_));
 sky130_fd_sc_hd__and3_1 _08994_ (.A(_00303_),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[38] ),
    .C(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__buf_2 _08995_ (.A(net25),
    .X(_03503_));
 sky130_fd_sc_hd__buf_2 _08996_ (.A(net26),
    .X(_03504_));
 sky130_fd_sc_hd__buf_2 _08997_ (.A(net12),
    .X(_03505_));
 sky130_fd_sc_hd__buf_2 _08998_ (.A(net13),
    .X(_03506_));
 sky130_fd_sc_hd__mux4_1 _08999_ (.A0(_03503_),
    .A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[36] ),
    .X(_03507_));
 sky130_fd_sc_hd__a31o_1 _09000_ (.A1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[37] ),
    .A2(_00307_),
    .A3(_03507_),
    .B1(_00309_),
    .X(_03508_));
 sky130_fd_sc_hd__a211oi_1 _09001_ (.A1(_03477_),
    .A2(_03492_),
    .B1(_03502_),
    .C1(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__a31oi_1 _09002_ (.A1(_03472_),
    .A2(_03476_),
    .A3(net3632),
    .B1(_03509_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[7] ));
 sky130_fd_sc_hd__inv_2 _09003_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[33] ),
    .Y(_03510_));
 sky130_fd_sc_hd__buf_2 _09004_ (.A(_01580_),
    .X(_03511_));
 sky130_fd_sc_hd__buf_2 _09005_ (.A(_01673_),
    .X(_03512_));
 sky130_fd_sc_hd__buf_2 _09006_ (.A(_01759_),
    .X(_03513_));
 sky130_fd_sc_hd__buf_2 _09007_ (.A(_01849_),
    .X(_03514_));
 sky130_fd_sc_hd__mux4_1 _09008_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ),
    .X(_03515_));
 sky130_fd_sc_hd__buf_2 _09009_ (.A(net11),
    .X(_03516_));
 sky130_fd_sc_hd__buf_2 _09010_ (.A(net18),
    .X(_03517_));
 sky130_fd_sc_hd__buf_2 _09011_ (.A(net19),
    .X(_03518_));
 sky130_fd_sc_hd__buf_2 _09012_ (.A(net20),
    .X(_03519_));
 sky130_fd_sc_hd__mux4_1 _09013_ (.A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ),
    .X(_03520_));
 sky130_fd_sc_hd__o21ai_1 _09014_ (.A1(_03510_),
    .A2(_03520_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[32] ),
    .Y(_03521_));
 sky130_fd_sc_hd__a21oi_1 _09015_ (.A1(_03510_),
    .A2(_03515_),
    .B1(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__nor2_1 _09016_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[32] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[33] ),
    .Y(_03523_));
 sky130_fd_sc_hd__buf_2 _09017_ (.A(_02226_),
    .X(_03524_));
 sky130_fd_sc_hd__buf_2 _09018_ (.A(_02320_),
    .X(_03525_));
 sky130_fd_sc_hd__buf_2 _09019_ (.A(_02408_),
    .X(_03526_));
 sky130_fd_sc_hd__buf_2 _09020_ (.A(_02491_),
    .X(_03527_));
 sky130_fd_sc_hd__mux4_1 _09021_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ),
    .X(_03528_));
 sky130_fd_sc_hd__a21o_1 _09022_ (.A1(_03523_),
    .A2(_03528_),
    .B1(net3764),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_4 _09023_ (.A(_00880_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_4 _09024_ (.A(_00972_),
    .X(_03531_));
 sky130_fd_sc_hd__buf_4 _09025_ (.A(_01311_),
    .X(_03532_));
 sky130_fd_sc_hd__buf_4 _09026_ (.A(_01395_),
    .X(_03533_));
 sky130_fd_sc_hd__mux4_1 _09027_ (.A0(_03530_),
    .A1(_03531_),
    .A2(_03532_),
    .A3(_03533_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ),
    .X(_03534_));
 sky130_fd_sc_hd__nor3_1 _09028_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[32] ),
    .B(_03510_),
    .C(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__buf_2 _09029_ (.A(_03484_),
    .X(_03536_));
 sky130_fd_sc_hd__buf_2 _09030_ (.A(_03486_),
    .X(_03537_));
 sky130_fd_sc_hd__buf_2 _09031_ (.A(_03488_),
    .X(_03538_));
 sky130_fd_sc_hd__buf_2 _09032_ (.A(_03490_),
    .X(_03539_));
 sky130_fd_sc_hd__mux4_1 _09033_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_4 _09034_ (.A(net25),
    .X(_03541_));
 sky130_fd_sc_hd__clkbuf_4 _09035_ (.A(net26),
    .X(_03542_));
 sky130_fd_sc_hd__clkbuf_4 _09036_ (.A(net12),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_4 _09037_ (.A(net13),
    .X(_03544_));
 sky130_fd_sc_hd__mux4_1 _09038_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ),
    .X(_03545_));
 sky130_fd_sc_hd__buf_2 _09039_ (.A(net14),
    .X(_03546_));
 sky130_fd_sc_hd__buf_2 _09040_ (.A(net15),
    .X(_03547_));
 sky130_fd_sc_hd__buf_2 _09041_ (.A(net16),
    .X(_03548_));
 sky130_fd_sc_hd__buf_2 _09042_ (.A(net17),
    .X(_03549_));
 sky130_fd_sc_hd__mux4_1 _09043_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ),
    .X(_03550_));
 sky130_fd_sc_hd__and3b_1 _09044_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[32] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[33] ),
    .C(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__a31o_1 _09045_ (.A1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[32] ),
    .A2(_03510_),
    .A3(_03545_),
    .B1(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__inv_2 _09046_ (.A(net3764),
    .Y(_03553_));
 sky130_fd_sc_hd__a211o_1 _09047_ (.A1(_03523_),
    .A2(_03540_),
    .B1(_03552_),
    .C1(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__o31a_1 _09048_ (.A1(_03522_),
    .A2(_03529_),
    .A3(_03535_),
    .B1(_03554_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[6] ));
 sky130_fd_sc_hd__inv_2 _09049_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[28] ),
    .Y(_03555_));
 sky130_fd_sc_hd__mux4_1 _09050_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ),
    .X(_03556_));
 sky130_fd_sc_hd__mux4_1 _09051_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ),
    .X(_03557_));
 sky130_fd_sc_hd__o21ai_1 _09052_ (.A1(_03555_),
    .A2(_03557_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[27] ),
    .Y(_03558_));
 sky130_fd_sc_hd__a21o_1 _09053_ (.A1(_03555_),
    .A2(_03556_),
    .B1(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__mux4_1 _09054_ (.A0(_00880_),
    .A1(_00972_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ),
    .X(_03560_));
 sky130_fd_sc_hd__or3_1 _09055_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[27] ),
    .B(_03555_),
    .C(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__nor2_1 _09056_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[27] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[28] ),
    .Y(_03562_));
 sky130_fd_sc_hd__mux4_1 _09057_ (.A0(_03478_),
    .A1(_03479_),
    .A2(_03480_),
    .A3(_03481_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ),
    .X(_03563_));
 sky130_fd_sc_hd__a21oi_1 _09058_ (.A1(_03562_),
    .A2(_03563_),
    .B1(net3494),
    .Y(_03564_));
 sky130_fd_sc_hd__mux4_1 _09059_ (.A0(_03485_),
    .A1(_03487_),
    .A2(_03489_),
    .A3(_03491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ),
    .X(_03565_));
 sky130_fd_sc_hd__mux4_1 _09060_ (.A0(_03494_),
    .A1(_03496_),
    .A2(_03498_),
    .A3(_03500_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ),
    .X(_03566_));
 sky130_fd_sc_hd__and3b_1 _09061_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[27] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[28] ),
    .C(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__mux4_1 _09062_ (.A0(_03503_),
    .A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ),
    .X(_03568_));
 sky130_fd_sc_hd__inv_2 _09063_ (.A(net3494),
    .Y(_03569_));
 sky130_fd_sc_hd__a31o_1 _09064_ (.A1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[27] ),
    .A2(_03555_),
    .A3(_03568_),
    .B1(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__a211oi_1 _09065_ (.A1(_03562_),
    .A2(_03565_),
    .B1(_03567_),
    .C1(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__a31oi_1 _09066_ (.A1(_03559_),
    .A2(_03561_),
    .A3(_03564_),
    .B1(_03571_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[5] ));
 sky130_fd_sc_hd__mux4_1 _09067_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ),
    .X(_03572_));
 sky130_fd_sc_hd__mux4_1 _09068_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ),
    .X(_03573_));
 sky130_fd_sc_hd__nor2_1 _09069_ (.A(_00274_),
    .B(_03573_),
    .Y(_03574_));
 sky130_fd_sc_hd__inv_2 _09070_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ),
    .Y(_03575_));
 sky130_fd_sc_hd__a211o_1 _09071_ (.A1(_00274_),
    .A2(_03572_),
    .B1(_03574_),
    .C1(_03575_),
    .X(_03576_));
 sky130_fd_sc_hd__mux4_1 _09072_ (.A0(_00880_),
    .A1(_00972_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ),
    .X(_03577_));
 sky130_fd_sc_hd__or3_1 _09073_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ),
    .B(_00274_),
    .C(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__nor2_1 _09074_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[23] ),
    .Y(_03579_));
 sky130_fd_sc_hd__mux4_1 _09075_ (.A0(_03478_),
    .A1(_03479_),
    .A2(_03480_),
    .A3(_03481_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ),
    .X(_03580_));
 sky130_fd_sc_hd__a21oi_1 _09076_ (.A1(_03579_),
    .A2(_03580_),
    .B1(net3390),
    .Y(_03581_));
 sky130_fd_sc_hd__mux4_1 _09077_ (.A0(net25),
    .A1(net26),
    .A2(net12),
    .A3(net13),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ),
    .X(_03582_));
 sky130_fd_sc_hd__or3b_1 _09078_ (.A(_03575_),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[23] ),
    .C_N(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__mux4_1 _09079_ (.A0(net21),
    .A1(net22),
    .A2(net23),
    .A3(net24),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ),
    .X(_03584_));
 sky130_fd_sc_hd__mux4_1 _09080_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ),
    .X(_03585_));
 sky130_fd_sc_hd__nand2_1 _09081_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[23] ),
    .B(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__o2bb2a_1 _09082_ (.A1_N(_03579_),
    .A2_N(_03584_),
    .B1(_03586_),
    .B2(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ),
    .X(_03587_));
 sky130_fd_sc_hd__and3_1 _09083_ (.A(net3390),
    .B(_03583_),
    .C(_03587_),
    .X(_03588_));
 sky130_fd_sc_hd__a31oi_1 _09084_ (.A1(_03576_),
    .A2(_03578_),
    .A3(net3391),
    .B1(_03588_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[4] ));
 sky130_fd_sc_hd__nand3b_2 _09085_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .B(_01415_),
    .C(net1),
    .Y(_03589_));
 sky130_fd_sc_hd__or3_1 _09086_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_03590_));
 sky130_fd_sc_hd__or2_1 _09087_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_03590_),
    .X(_03591_));
 sky130_fd_sc_hd__o21a_2 _09088_ (.A1(_03589_),
    .A2(_03591_),
    .B1(_03013_),
    .X(_03592_));
 sky130_fd_sc_hd__mux2_1 _09089_ (.A0(_03344_),
    .A1(net3497),
    .S(_03592_),
    .X(_03593_));
 sky130_fd_sc_hd__clkbuf_1 _09090_ (.A(_03593_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__inv_2 _09091_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[18] ),
    .Y(_03594_));
 sky130_fd_sc_hd__mux4_1 _09092_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[16] ),
    .X(_03595_));
 sky130_fd_sc_hd__mux4_1 _09093_ (.A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[16] ),
    .X(_03596_));
 sky130_fd_sc_hd__o21ai_1 _09094_ (.A1(_03594_),
    .A2(_03596_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[17] ),
    .Y(_03597_));
 sky130_fd_sc_hd__a21oi_1 _09095_ (.A1(_03594_),
    .A2(_03595_),
    .B1(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__mux4_1 _09096_ (.A0(_03530_),
    .A1(_03531_),
    .A2(_03532_),
    .A3(_03533_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[16] ),
    .X(_03599_));
 sky130_fd_sc_hd__nor3_1 _09097_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[17] ),
    .B(_03594_),
    .C(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__nor2_1 _09098_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[17] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[18] ),
    .Y(_03601_));
 sky130_fd_sc_hd__mux4_1 _09099_ (.A0(_03478_),
    .A1(_03479_),
    .A2(_03480_),
    .A3(_03481_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[16] ),
    .X(_03602_));
 sky130_fd_sc_hd__a21o_1 _09100_ (.A1(_03601_),
    .A2(_03602_),
    .B1(net3725),
    .X(_03603_));
 sky130_fd_sc_hd__mux4_1 _09101_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[16] ),
    .X(_03604_));
 sky130_fd_sc_hd__mux4_1 _09102_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[16] ),
    .X(_03605_));
 sky130_fd_sc_hd__mux4_1 _09103_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[16] ),
    .X(_03606_));
 sky130_fd_sc_hd__and3b_1 _09104_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[17] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[18] ),
    .C(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__a31o_1 _09105_ (.A1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[17] ),
    .A2(_03594_),
    .A3(_03605_),
    .B1(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__inv_2 _09106_ (.A(net3725),
    .Y(_03609_));
 sky130_fd_sc_hd__a211o_1 _09107_ (.A1(_03601_),
    .A2(_03604_),
    .B1(_03608_),
    .C1(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__o31a_1 _09108_ (.A1(_03598_),
    .A2(_03600_),
    .A3(_03603_),
    .B1(_03610_),
    .X(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[3] ));
 sky130_fd_sc_hd__mux2_1 _09109_ (.A0(_03351_),
    .A1(net3327),
    .S(_03592_),
    .X(_03611_));
 sky130_fd_sc_hd__clkbuf_1 _09110_ (.A(_03611_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _09111_ (.A0(_03353_),
    .A1(net3381),
    .S(_03592_),
    .X(_03612_));
 sky130_fd_sc_hd__clkbuf_1 _09112_ (.A(_03612_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _09113_ (.A0(_03246_),
    .A1(net3512),
    .S(_03592_),
    .X(_03613_));
 sky130_fd_sc_hd__clkbuf_1 _09114_ (.A(_03613_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _09115_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_2 _09116_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ),
    .X(_03615_));
 sky130_fd_sc_hd__inv_2 _09117_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .Y(_03616_));
 sky130_fd_sc_hd__or4_1 _09118_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_03615_),
    .C(_03616_),
    .D(_03589_),
    .X(_03617_));
 sky130_fd_sc_hd__o21a_2 _09119_ (.A1(_03614_),
    .A2(_03617_),
    .B1(_03013_),
    .X(_03618_));
 sky130_fd_sc_hd__mux2_1 _09120_ (.A0(_03344_),
    .A1(net3574),
    .S(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__clkbuf_1 _09121_ (.A(_03619_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _09122_ (.A0(_03351_),
    .A1(net3434),
    .S(_03618_),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_1 _09123_ (.A(_03620_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _09124_ (.A0(_03353_),
    .A1(net3814),
    .S(_03618_),
    .X(_03621_));
 sky130_fd_sc_hd__clkbuf_1 _09125_ (.A(_03621_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__buf_4 _09126_ (.A(_00191_),
    .X(_03622_));
 sky130_fd_sc_hd__mux2_1 _09127_ (.A0(_03622_),
    .A1(net3614),
    .S(_03618_),
    .X(_03623_));
 sky130_fd_sc_hd__clkbuf_1 _09128_ (.A(_03623_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__and3b_2 _09129_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .B(_01415_),
    .C(net1),
    .X(_03624_));
 sky130_fd_sc_hd__nand2_1 _09130_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_03590_),
    .Y(_03625_));
 sky130_fd_sc_hd__and2_1 _09131_ (.A(_03591_),
    .B(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__inv_2 _09132_ (.A(_03614_),
    .Y(_03627_));
 sky130_fd_sc_hd__or3_1 _09133_ (.A(_03615_),
    .B(_03627_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_03628_));
 sky130_fd_sc_hd__nand2_1 _09134_ (.A(_00170_),
    .B(_03591_),
    .Y(_03629_));
 sky130_fd_sc_hd__nor2_1 _09135_ (.A(_03628_),
    .B(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__inv_2 _09136_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .Y(_03631_));
 sky130_fd_sc_hd__and3b_2 _09137_ (.A_N(_03628_),
    .B(_03631_),
    .C(_03624_),
    .X(_03632_));
 sky130_fd_sc_hd__inv_2 _09138_ (.A(_03632_),
    .Y(_03633_));
 sky130_fd_sc_hd__a32o_1 _09139_ (.A1(_03624_),
    .A2(_03626_),
    .A3(_03630_),
    .B1(_03633_),
    .B2(net3815),
    .X(_03634_));
 sky130_fd_sc_hd__a21o_1 _09140_ (.A1(_02044_),
    .A2(_03634_),
    .B1(_00210_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__clkinv_2 _09141_ (.A(net3569),
    .Y(_03635_));
 sky130_fd_sc_hd__nand2_1 _09142_ (.A(_01446_),
    .B(_03591_),
    .Y(_03636_));
 sky130_fd_sc_hd__mux2_1 _09143_ (.A0(_03635_),
    .A1(_03636_),
    .S(_03632_),
    .X(_03637_));
 sky130_fd_sc_hd__o21ai_1 _09144_ (.A1(_03408_),
    .A2(_03637_),
    .B1(_03379_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__and2_1 _09145_ (.A(_00187_),
    .B(_03591_),
    .X(_03638_));
 sky130_fd_sc_hd__mux2_1 _09146_ (.A0(net3816),
    .A1(_03638_),
    .S(_03632_),
    .X(_03639_));
 sky130_fd_sc_hd__a21o_1 _09147_ (.A1(_02044_),
    .A2(_03639_),
    .B1(_00262_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__clkinv_2 _09148_ (.A(net3445),
    .Y(_03640_));
 sky130_fd_sc_hd__nand2_1 _09149_ (.A(_01452_),
    .B(_03591_),
    .Y(_03641_));
 sky130_fd_sc_hd__mux2_1 _09150_ (.A0(_03640_),
    .A1(_03641_),
    .S(_03632_),
    .X(_03642_));
 sky130_fd_sc_hd__o21ai_1 _09151_ (.A1(_03408_),
    .A2(_03642_),
    .B1(_03322_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _09152_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(_03589_),
    .Y(_03643_));
 sky130_fd_sc_hd__and3b_2 _09153_ (.A_N(_03615_),
    .B(_03614_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(_03644_));
 sky130_fd_sc_hd__a21oi_4 _09154_ (.A1(_03643_),
    .A2(_03644_),
    .B1(_02686_),
    .Y(_03645_));
 sky130_fd_sc_hd__mux2_1 _09155_ (.A0(_03344_),
    .A1(net3476),
    .S(_03645_),
    .X(_03646_));
 sky130_fd_sc_hd__clkbuf_1 _09156_ (.A(_03646_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _09157_ (.A0(_03351_),
    .A1(net3622),
    .S(_03645_),
    .X(_03647_));
 sky130_fd_sc_hd__clkbuf_1 _09158_ (.A(_03647_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _09159_ (.A0(_03353_),
    .A1(net3561),
    .S(_03645_),
    .X(_03648_));
 sky130_fd_sc_hd__clkbuf_1 _09160_ (.A(_03648_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__inv_2 _09161_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[13] ),
    .Y(_03649_));
 sky130_fd_sc_hd__mux4_1 _09162_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ),
    .X(_03650_));
 sky130_fd_sc_hd__mux4_1 _09163_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ),
    .X(_03651_));
 sky130_fd_sc_hd__nor2_1 _09164_ (.A(_03649_),
    .B(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__a211o_1 _09165_ (.A1(_03649_),
    .A2(_03650_),
    .B1(_03652_),
    .C1(_00242_),
    .X(_03653_));
 sky130_fd_sc_hd__mux4_1 _09166_ (.A0(_00880_),
    .A1(_00972_),
    .A2(_01311_),
    .A3(_01395_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ),
    .X(_03654_));
 sky130_fd_sc_hd__or3_1 _09167_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[12] ),
    .B(_03649_),
    .C(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__nor2_1 _09168_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[12] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[13] ),
    .Y(_03656_));
 sky130_fd_sc_hd__mux4_1 _09169_ (.A0(_03478_),
    .A1(_03479_),
    .A2(_03480_),
    .A3(_03481_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ),
    .X(_03657_));
 sky130_fd_sc_hd__a21oi_1 _09170_ (.A1(_03656_),
    .A2(_03657_),
    .B1(net3663),
    .Y(_03658_));
 sky130_fd_sc_hd__mux4_1 _09171_ (.A0(_03485_),
    .A1(_03487_),
    .A2(_03489_),
    .A3(_03491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ),
    .X(_03659_));
 sky130_fd_sc_hd__mux4_1 _09172_ (.A0(_03494_),
    .A1(_03496_),
    .A2(_03498_),
    .A3(_03500_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ),
    .X(_03660_));
 sky130_fd_sc_hd__and3_1 _09173_ (.A(_00242_),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[13] ),
    .C(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__mux4_1 _09174_ (.A0(_03503_),
    .A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ),
    .X(_03662_));
 sky130_fd_sc_hd__a31o_1 _09175_ (.A1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[12] ),
    .A2(_03649_),
    .A3(_03662_),
    .B1(_00247_),
    .X(_03663_));
 sky130_fd_sc_hd__a211oi_1 _09176_ (.A1(_03656_),
    .A2(_03659_),
    .B1(_03661_),
    .C1(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__a31oi_1 _09177_ (.A1(_03653_),
    .A2(_03655_),
    .A3(net3664),
    .B1(_03664_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[2] ));
 sky130_fd_sc_hd__mux2_1 _09178_ (.A0(_03622_),
    .A1(net3563),
    .S(_03645_),
    .X(_03665_));
 sky130_fd_sc_hd__clkbuf_1 _09179_ (.A(_03665_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__clkbuf_4 _09180_ (.A(_00195_),
    .X(_03666_));
 sky130_fd_sc_hd__and4_1 _09181_ (.A(_03615_),
    .B(_03627_),
    .C(_03616_),
    .D(_03643_),
    .X(_03667_));
 sky130_fd_sc_hd__clkbuf_2 _09182_ (.A(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__nand2_1 _09183_ (.A(_03629_),
    .B(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__or2_1 _09184_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .B(_03668_),
    .X(_03670_));
 sky130_fd_sc_hd__a31o_1 _09185_ (.A1(_03666_),
    .A2(_03669_),
    .A3(_03670_),
    .B1(_03316_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _09186_ (.A(_03636_),
    .B(_03668_),
    .Y(_03671_));
 sky130_fd_sc_hd__or2_1 _09187_ (.A(net3217),
    .B(_03668_),
    .X(_03672_));
 sky130_fd_sc_hd__a31o_1 _09188_ (.A1(_03666_),
    .A2(_03671_),
    .A3(_03672_),
    .B1(_03050_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__or2b_1 _09189_ (.A(_03638_),
    .B_N(_03668_),
    .X(_03673_));
 sky130_fd_sc_hd__or2_1 _09190_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .B(_03668_),
    .X(_03674_));
 sky130_fd_sc_hd__a31o_1 _09191_ (.A1(_03666_),
    .A2(_03673_),
    .A3(_03674_),
    .B1(_01851_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _09192_ (.A(net3991),
    .B(_03668_),
    .Y(_03675_));
 sky130_fd_sc_hd__a211o_1 _09193_ (.A1(_03641_),
    .A2(_03668_),
    .B1(_03675_),
    .C1(_02868_),
    .X(_03676_));
 sky130_fd_sc_hd__nand2_1 _09194_ (.A(_03166_),
    .B(_03676_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _09195_ (.A1(_03615_),
    .A2(_03627_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .A4(_03643_),
    .B1(_00249_),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_1 _09196_ (.A0(net4045),
    .A1(_03169_),
    .S(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_1 _09197_ (.A(_03678_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(net4199),
    .A1(_03172_),
    .S(_03677_),
    .X(_03679_));
 sky130_fd_sc_hd__clkbuf_1 _09199_ (.A(_03679_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(net4005),
    .A1(_03174_),
    .S(_03677_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_1 _09201_ (.A(_03680_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _09202_ (.A0(net3493),
    .A1(_00527_),
    .S(_03677_),
    .X(_03681_));
 sky130_fd_sc_hd__clkbuf_1 _09203_ (.A(_03681_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_2 _09204_ (.A(_03615_),
    .B(_03614_),
    .C(_03616_),
    .D(_03643_),
    .X(_03682_));
 sky130_fd_sc_hd__or2_1 _09205_ (.A(net4132),
    .B(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__nand2_1 _09206_ (.A(_03629_),
    .B(_03682_),
    .Y(_03684_));
 sky130_fd_sc_hd__a31o_1 _09207_ (.A1(_03666_),
    .A2(_03683_),
    .A3(_03684_),
    .B1(_03316_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _09208_ (.A0(_01161_),
    .A1(_03636_),
    .S(_03682_),
    .X(_03685_));
 sky130_fd_sc_hd__o21ai_1 _09209_ (.A1(_03408_),
    .A2(_03685_),
    .B1(_03379_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _09210_ (.A0(net4173),
    .A1(_03638_),
    .S(_03682_),
    .X(_03686_));
 sky130_fd_sc_hd__a21o_1 _09211_ (.A1(_02044_),
    .A2(_03686_),
    .B1(_00262_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _09212_ (.A0(_01153_),
    .A1(_03641_),
    .S(_03682_),
    .X(_03687_));
 sky130_fd_sc_hd__o21ai_1 _09213_ (.A1(_03408_),
    .A2(_03687_),
    .B1(_03322_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _09214_ (.A1(_03615_),
    .A2(_03614_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .A4(_03643_),
    .B1(_00249_),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _09215_ (.A0(net4202),
    .A1(_03169_),
    .S(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__clkbuf_1 _09216_ (.A(_03689_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux4_1 _09217_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ),
    .X(_03690_));
 sky130_fd_sc_hd__mux4_1 _09218_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ),
    .X(_03691_));
 sky130_fd_sc_hd__o21ai_1 _09219_ (.A1(_00230_),
    .A2(_03691_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ),
    .Y(_03692_));
 sky130_fd_sc_hd__a21o_1 _09220_ (.A1(_00230_),
    .A2(_03690_),
    .B1(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__nor2_1 _09221_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[8] ),
    .Y(_03694_));
 sky130_fd_sc_hd__mux4_1 _09222_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ),
    .X(_03695_));
 sky130_fd_sc_hd__a21oi_1 _09223_ (.A1(_03694_),
    .A2(_03695_),
    .B1(net3488),
    .Y(_03696_));
 sky130_fd_sc_hd__buf_4 _09224_ (.A(_00879_),
    .X(_03697_));
 sky130_fd_sc_hd__clkbuf_4 _09225_ (.A(_00972_),
    .X(_03698_));
 sky130_fd_sc_hd__mux4_1 _09226_ (.A0(_03697_),
    .A1(_03698_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ),
    .X(_03699_));
 sky130_fd_sc_hd__or3_1 _09227_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ),
    .B(_00230_),
    .C(_03699_),
    .X(_03700_));
 sky130_fd_sc_hd__mux4_1 _09228_ (.A0(_03485_),
    .A1(_03487_),
    .A2(_03489_),
    .A3(_03491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ),
    .X(_03701_));
 sky130_fd_sc_hd__mux4_1 _09229_ (.A0(_03494_),
    .A1(_03496_),
    .A2(_03498_),
    .A3(_03500_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ),
    .X(_03702_));
 sky130_fd_sc_hd__and3b_1 _09230_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[8] ),
    .C(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__mux4_1 _09231_ (.A0(_03503_),
    .A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ),
    .X(_03704_));
 sky130_fd_sc_hd__inv_2 _09232_ (.A(net3488),
    .Y(_03705_));
 sky130_fd_sc_hd__a31o_1 _09233_ (.A1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ),
    .A2(_00230_),
    .A3(_03704_),
    .B1(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__a211oi_1 _09234_ (.A1(_03694_),
    .A2(_03701_),
    .B1(_03703_),
    .C1(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__a31oi_1 _09235_ (.A1(_03693_),
    .A2(net3489),
    .A3(_03700_),
    .B1(_03707_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[1] ));
 sky130_fd_sc_hd__mux2_1 _09236_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .A1(_03172_),
    .S(_03688_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_1 _09237_ (.A(_03708_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _09238_ (.A0(net3763),
    .A1(_03174_),
    .S(_03688_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_1 _09239_ (.A(_03709_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _09240_ (.A0(net3897),
    .A1(_00527_),
    .S(_03688_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_1 _09241_ (.A(_03710_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__o31a_2 _09242_ (.A1(_03631_),
    .A2(_03589_),
    .A3(_03590_),
    .B1(_02847_),
    .X(_03711_));
 sky130_fd_sc_hd__mux2_1 _09243_ (.A0(_03344_),
    .A1(net3957),
    .S(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__clkbuf_1 _09244_ (.A(_03712_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _09245_ (.A0(_03351_),
    .A1(net3148),
    .S(_03711_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_1 _09246_ (.A(_03713_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _09247_ (.A0(_03353_),
    .A1(net3770),
    .S(_03711_),
    .X(_03714_));
 sky130_fd_sc_hd__clkbuf_1 _09248_ (.A(_03714_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _09249_ (.A0(_03622_),
    .A1(net3829),
    .S(_03711_),
    .X(_03715_));
 sky130_fd_sc_hd__clkbuf_1 _09250_ (.A(_03715_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _09251_ (.A(_03589_),
    .B(_03626_),
    .X(_03716_));
 sky130_fd_sc_hd__o41a_2 _09252_ (.A1(_03615_),
    .A2(_03614_),
    .A3(_03616_),
    .A4(_03716_),
    .B1(_00407_),
    .X(_03717_));
 sky130_fd_sc_hd__mux2_1 _09253_ (.A0(_03344_),
    .A1(net3834),
    .S(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_1 _09254_ (.A(_03718_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _09255_ (.A0(_03351_),
    .A1(net3171),
    .S(_03717_),
    .X(_03719_));
 sky130_fd_sc_hd__clkbuf_1 _09256_ (.A(_03719_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _09257_ (.A0(_03353_),
    .A1(net3742),
    .S(_03717_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_1 _09258_ (.A(_03720_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _09259_ (.A0(_03622_),
    .A1(net3516),
    .S(_03717_),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_1 _09260_ (.A(_03721_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _09261_ (.A(_03628_),
    .B(_03716_),
    .Y(_03722_));
 sky130_fd_sc_hd__or2_1 _09262_ (.A(net4153),
    .B(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__nand2_1 _09263_ (.A(_03629_),
    .B(_03722_),
    .Y(_03724_));
 sky130_fd_sc_hd__a31o_1 _09264_ (.A1(_03666_),
    .A2(_03723_),
    .A3(_03724_),
    .B1(_03316_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__nand2_1 _09265_ (.A(_03636_),
    .B(_03722_),
    .Y(_03725_));
 sky130_fd_sc_hd__or2_1 _09266_ (.A(net4046),
    .B(_03722_),
    .X(_03726_));
 sky130_fd_sc_hd__a31o_1 _09267_ (.A1(_03666_),
    .A2(_03725_),
    .A3(_03726_),
    .B1(_03050_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__mux2_1 _09268_ (.A0(net3140),
    .A1(_03638_),
    .S(_03722_),
    .X(_03727_));
 sky130_fd_sc_hd__a21o_1 _09269_ (.A1(_02044_),
    .A2(_03727_),
    .B1(_00262_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__inv_2 _09270_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[3] ),
    .Y(_03728_));
 sky130_fd_sc_hd__mux4_1 _09271_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[1] ),
    .X(_03729_));
 sky130_fd_sc_hd__mux4_1 _09272_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[1] ),
    .X(_03730_));
 sky130_fd_sc_hd__o21ai_1 _09273_ (.A1(_03728_),
    .A2(_03730_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[2] ),
    .Y(_03731_));
 sky130_fd_sc_hd__a21o_1 _09274_ (.A1(_03728_),
    .A2(_03729_),
    .B1(_03731_),
    .X(_03732_));
 sky130_fd_sc_hd__mux4_1 _09275_ (.A0(_00880_),
    .A1(_00972_),
    .A2(_01311_),
    .A3(_01395_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[1] ),
    .X(_03733_));
 sky130_fd_sc_hd__or3_1 _09276_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[2] ),
    .B(_03728_),
    .C(_03733_),
    .X(_03734_));
 sky130_fd_sc_hd__nor2_1 _09277_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[2] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[3] ),
    .Y(_03735_));
 sky130_fd_sc_hd__mux4_1 _09278_ (.A0(_03478_),
    .A1(_03479_),
    .A2(_03480_),
    .A3(_03481_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[1] ),
    .X(_03736_));
 sky130_fd_sc_hd__a21oi_1 _09279_ (.A1(_03735_),
    .A2(_03736_),
    .B1(net3415),
    .Y(_03737_));
 sky130_fd_sc_hd__mux4_1 _09280_ (.A0(_03485_),
    .A1(_03487_),
    .A2(_03489_),
    .A3(_03491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[1] ),
    .X(_03738_));
 sky130_fd_sc_hd__mux4_1 _09281_ (.A0(_03494_),
    .A1(_03496_),
    .A2(_03498_),
    .A3(_03500_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[1] ),
    .X(_03739_));
 sky130_fd_sc_hd__and3b_1 _09282_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[2] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[3] ),
    .C(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__mux4_1 _09283_ (.A0(_03503_),
    .A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[1] ),
    .X(_03741_));
 sky130_fd_sc_hd__inv_2 _09284_ (.A(net3415),
    .Y(_03742_));
 sky130_fd_sc_hd__a31o_1 _09285_ (.A1(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[2] ),
    .A2(_03728_),
    .A3(_03741_),
    .B1(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__a211oi_1 _09286_ (.A1(_03735_),
    .A2(_03738_),
    .B1(_03740_),
    .C1(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__a31oi_1 _09287_ (.A1(_03732_),
    .A2(_03734_),
    .A3(net3416),
    .B1(_03744_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[0] ));
 sky130_fd_sc_hd__nor2_1 _09288_ (.A(net4105),
    .B(_03722_),
    .Y(_03745_));
 sky130_fd_sc_hd__a211o_1 _09289_ (.A1(_03641_),
    .A2(_03722_),
    .B1(_03745_),
    .C1(_02868_),
    .X(_03746_));
 sky130_fd_sc_hd__nand2_1 _09290_ (.A(_03166_),
    .B(_03746_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3b_1 _09291_ (.A_N(_03626_),
    .B(_03644_),
    .C(_03624_),
    .X(_03747_));
 sky130_fd_sc_hd__a31oi_4 _09292_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .A2(_03624_),
    .A3(_03644_),
    .B1(_02637_),
    .Y(_03748_));
 sky130_fd_sc_hd__a221o_1 _09293_ (.A1(_00288_),
    .A2(_03747_),
    .B1(_03748_),
    .B2(net3322),
    .C1(_00209_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _09294_ (.A1(_00293_),
    .A2(_03747_),
    .B1(_03748_),
    .B2(net3228),
    .C1(_02872_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _09295_ (.A1(_00295_),
    .A2(_03747_),
    .B1(_03748_),
    .B2(net3314),
    .C1(_00221_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__and2_1 _09296_ (.A(_01858_),
    .B(_01141_),
    .X(_03749_));
 sky130_fd_sc_hd__a22o_1 _09297_ (.A1(_01165_),
    .A2(_01218_),
    .B1(_01220_),
    .B2(_01224_),
    .X(_03750_));
 sky130_fd_sc_hd__and2_1 _09298_ (.A(_01578_),
    .B(_03750_),
    .X(_03751_));
 sky130_fd_sc_hd__mux2_1 _09299_ (.A0(_03749_),
    .A1(_03751_),
    .S(_01863_),
    .X(_03752_));
 sky130_fd_sc_hd__clkbuf_1 _09300_ (.A(_03752_),
    .X(_00000_));
 sky130_fd_sc_hd__inv_2 _09301_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ),
    .Y(_03753_));
 sky130_fd_sc_hd__mux4_1 _09302_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ),
    .X(_03754_));
 sky130_fd_sc_hd__mux4_1 _09303_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ),
    .X(_03755_));
 sky130_fd_sc_hd__o21ai_1 _09304_ (.A1(_03753_),
    .A2(_03755_),
    .B1(net3842),
    .Y(_03756_));
 sky130_fd_sc_hd__a21o_1 _09305_ (.A1(_03753_),
    .A2(_03754_),
    .B1(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_4 _09306_ (.A(_01227_),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_4 _09307_ (.A(_01056_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_4 _09308_ (.A(_00784_),
    .X(_03760_));
 sky130_fd_sc_hd__clkbuf_4 _09309_ (.A(_01143_),
    .X(_03761_));
 sky130_fd_sc_hd__mux4_1 _09310_ (.A0(_03758_),
    .A1(_03759_),
    .A2(_03760_),
    .A3(_03761_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[35] ),
    .X(_03762_));
 sky130_fd_sc_hd__inv_2 _09311_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[39] ),
    .Y(_03763_));
 sky130_fd_sc_hd__o31a_1 _09312_ (.A1(net3842),
    .A2(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ),
    .A3(_03762_),
    .B1(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__mux4_1 _09313_ (.A0(_03697_),
    .A1(_03698_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ),
    .X(_03765_));
 sky130_fd_sc_hd__or3_1 _09314_ (.A(net3842),
    .B(_03753_),
    .C(_03765_),
    .X(_03766_));
 sky130_fd_sc_hd__mux4_1 _09315_ (.A0(_03484_),
    .A1(_03486_),
    .A2(_03488_),
    .A3(_03490_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ),
    .X(_03767_));
 sky130_fd_sc_hd__inv_2 _09316_ (.A(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__mux4_1 _09317_ (.A0(_03503_),
    .A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ),
    .X(_03769_));
 sky130_fd_sc_hd__mux4_1 _09318_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ),
    .X(_03770_));
 sky130_fd_sc_hd__and3b_1 _09319_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[37] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ),
    .C(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__a31oi_1 _09320_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[37] ),
    .A2(_03753_),
    .A3(_03769_),
    .B1(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__o311a_1 _09321_ (.A1(net3842),
    .A2(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ),
    .A3(_03768_),
    .B1(_03772_),
    .C1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[39] ),
    .X(_03773_));
 sky130_fd_sc_hd__a31oi_1 _09322_ (.A1(_03757_),
    .A2(_03764_),
    .A3(net3843),
    .B1(_03773_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[7] ));
 sky130_fd_sc_hd__inv_2 _09323_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[33] ),
    .Y(_03774_));
 sky130_fd_sc_hd__mux4_1 _09324_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ),
    .X(_03775_));
 sky130_fd_sc_hd__mux4_1 _09325_ (.A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ),
    .X(_03776_));
 sky130_fd_sc_hd__o21ai_1 _09326_ (.A1(_03774_),
    .A2(_03776_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[32] ),
    .Y(_03777_));
 sky130_fd_sc_hd__a21oi_1 _09327_ (.A1(_03774_),
    .A2(_03775_),
    .B1(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__nor2_1 _09328_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[32] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[33] ),
    .Y(_03779_));
 sky130_fd_sc_hd__clkbuf_4 _09329_ (.A(_00785_),
    .X(_03780_));
 sky130_fd_sc_hd__clkbuf_4 _09330_ (.A(_01144_),
    .X(_03781_));
 sky130_fd_sc_hd__clkbuf_4 _09331_ (.A(_01228_),
    .X(_03782_));
 sky130_fd_sc_hd__clkbuf_4 _09332_ (.A(_01057_),
    .X(_03783_));
 sky130_fd_sc_hd__mux4_1 _09333_ (.A0(_03780_),
    .A1(_03781_),
    .A2(_03782_),
    .A3(_03783_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ),
    .S1(_00402_),
    .X(_03784_));
 sky130_fd_sc_hd__and2_1 _09334_ (.A(_03779_),
    .B(_03784_),
    .X(_03785_));
 sky130_fd_sc_hd__buf_4 _09335_ (.A(_01311_),
    .X(_03786_));
 sky130_fd_sc_hd__buf_4 _09336_ (.A(_01395_),
    .X(_03787_));
 sky130_fd_sc_hd__mux4_1 _09337_ (.A0(_03530_),
    .A1(_03531_),
    .A2(_03786_),
    .A3(_03787_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ),
    .X(_03788_));
 sky130_fd_sc_hd__nor3_1 _09338_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[32] ),
    .B(_03774_),
    .C(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__mux4_1 _09339_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ),
    .X(_03790_));
 sky130_fd_sc_hd__mux4_1 _09340_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ),
    .X(_03791_));
 sky130_fd_sc_hd__and3b_1 _09341_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[32] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[33] ),
    .C(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__mux4_1 _09342_ (.A0(_03503_),
    .A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ),
    .X(_03793_));
 sky130_fd_sc_hd__inv_2 _09343_ (.A(net3317),
    .Y(_03794_));
 sky130_fd_sc_hd__a31o_1 _09344_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[32] ),
    .A2(_03774_),
    .A3(_03793_),
    .B1(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__a211o_1 _09345_ (.A1(_03779_),
    .A2(_03790_),
    .B1(_03792_),
    .C1(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__o41a_1 _09346_ (.A1(net3317),
    .A2(_03778_),
    .A3(_03785_),
    .A4(_03789_),
    .B1(_03796_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[6] ));
 sky130_fd_sc_hd__mux4_1 _09347_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ),
    .X(_03797_));
 sky130_fd_sc_hd__mux4_1 _09348_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ),
    .X(_03798_));
 sky130_fd_sc_hd__nor2_1 _09349_ (.A(_00397_),
    .B(_03798_),
    .Y(_03799_));
 sky130_fd_sc_hd__a211o_1 _09350_ (.A1(_00397_),
    .A2(_03797_),
    .B1(_03799_),
    .C1(_00395_),
    .X(_03800_));
 sky130_fd_sc_hd__mux4_1 _09351_ (.A0(_03760_),
    .A1(_03761_),
    .A2(_03758_),
    .A3(_03759_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ),
    .S1(_00390_),
    .X(_03801_));
 sky130_fd_sc_hd__or3_1 _09352_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[27] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[28] ),
    .C(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__mux4_1 _09353_ (.A0(_03697_),
    .A1(_03698_),
    .A2(_03786_),
    .A3(_03787_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ),
    .X(_03803_));
 sky130_fd_sc_hd__o31a_1 _09354_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[27] ),
    .A2(_00397_),
    .A3(_03803_),
    .B1(_00400_),
    .X(_03804_));
 sky130_fd_sc_hd__mux4_1 _09355_ (.A0(_03485_),
    .A1(_03487_),
    .A2(_03489_),
    .A3(_03491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ),
    .X(_03805_));
 sky130_fd_sc_hd__clkbuf_4 _09356_ (.A(net25),
    .X(_03806_));
 sky130_fd_sc_hd__clkbuf_4 _09357_ (.A(net26),
    .X(_03807_));
 sky130_fd_sc_hd__clkbuf_4 _09358_ (.A(net12),
    .X(_03808_));
 sky130_fd_sc_hd__clkbuf_4 _09359_ (.A(net13),
    .X(_03809_));
 sky130_fd_sc_hd__mux4_1 _09360_ (.A0(_03806_),
    .A1(_03807_),
    .A2(_03808_),
    .A3(_03809_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ),
    .X(_03810_));
 sky130_fd_sc_hd__mux4_1 _09361_ (.A0(_03493_),
    .A1(_03495_),
    .A2(_03497_),
    .A3(_03499_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ),
    .X(_03811_));
 sky130_fd_sc_hd__and3_1 _09362_ (.A(_00395_),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[28] ),
    .C(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__a31o_1 _09363_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[27] ),
    .A2(_00397_),
    .A3(_03810_),
    .B1(_03812_),
    .X(_03813_));
 sky130_fd_sc_hd__a311oi_1 _09364_ (.A1(_00395_),
    .A2(_00397_),
    .A3(_03805_),
    .B1(_03813_),
    .C1(_00400_),
    .Y(_03814_));
 sky130_fd_sc_hd__a31oi_1 _09365_ (.A1(_03800_),
    .A2(_03802_),
    .A3(_03804_),
    .B1(net3576),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[5] ));
 sky130_fd_sc_hd__mux4_1 _09366_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_4 _09367_ (.A(net11),
    .X(_03816_));
 sky130_fd_sc_hd__buf_2 _09368_ (.A(net18),
    .X(_03817_));
 sky130_fd_sc_hd__clkbuf_4 _09369_ (.A(net19),
    .X(_03818_));
 sky130_fd_sc_hd__buf_2 _09370_ (.A(net20),
    .X(_03819_));
 sky130_fd_sc_hd__mux4_1 _09371_ (.A0(_03816_),
    .A1(_03817_),
    .A2(_03818_),
    .A3(_03819_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ),
    .X(_03820_));
 sky130_fd_sc_hd__nor2_1 _09372_ (.A(_00385_),
    .B(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__a211o_1 _09373_ (.A1(_00385_),
    .A2(_03815_),
    .B1(_03821_),
    .C1(_00383_),
    .X(_03822_));
 sky130_fd_sc_hd__mux4_1 _09374_ (.A0(_03760_),
    .A1(_03761_),
    .A2(_03758_),
    .A3(_03759_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ),
    .S1(_00377_),
    .X(_03823_));
 sky130_fd_sc_hd__o31a_1 _09375_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[22] ),
    .A2(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[23] ),
    .A3(_03823_),
    .B1(_00387_),
    .X(_03824_));
 sky130_fd_sc_hd__mux4_1 _09376_ (.A0(_03697_),
    .A1(_03698_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ),
    .X(_03825_));
 sky130_fd_sc_hd__or3_1 _09377_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[22] ),
    .B(_00385_),
    .C(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__mux4_1 _09378_ (.A0(_03485_),
    .A1(_03487_),
    .A2(_03489_),
    .A3(_03491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ),
    .X(_03827_));
 sky130_fd_sc_hd__mux4_1 _09379_ (.A0(_03806_),
    .A1(_03807_),
    .A2(_03808_),
    .A3(_03809_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ),
    .X(_03828_));
 sky130_fd_sc_hd__mux4_1 _09380_ (.A0(_03493_),
    .A1(_03495_),
    .A2(_03497_),
    .A3(_03499_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ),
    .X(_03829_));
 sky130_fd_sc_hd__and3_1 _09381_ (.A(_00383_),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[23] ),
    .C(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__a31o_1 _09382_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[22] ),
    .A2(_00385_),
    .A3(_03828_),
    .B1(_03830_),
    .X(_03831_));
 sky130_fd_sc_hd__a311oi_1 _09383_ (.A1(_00383_),
    .A2(_00385_),
    .A3(_03827_),
    .B1(_03831_),
    .C1(_00387_),
    .Y(_03832_));
 sky130_fd_sc_hd__a31oi_1 _09384_ (.A1(_03822_),
    .A2(_03824_),
    .A3(_03826_),
    .B1(net3701),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[4] ));
 sky130_fd_sc_hd__inv_2 _09385_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[18] ),
    .Y(_03833_));
 sky130_fd_sc_hd__mux4_1 _09386_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ),
    .X(_03834_));
 sky130_fd_sc_hd__mux4_1 _09387_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ),
    .X(_03835_));
 sky130_fd_sc_hd__o21ai_1 _09388_ (.A1(_03833_),
    .A2(_03835_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[17] ),
    .Y(_03836_));
 sky130_fd_sc_hd__a21o_1 _09389_ (.A1(_03833_),
    .A2(_03834_),
    .B1(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__mux4_1 _09390_ (.A0(_00784_),
    .A1(_01143_),
    .A2(_01227_),
    .A3(_01056_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ),
    .S1(_00365_),
    .X(_03838_));
 sky130_fd_sc_hd__or3_1 _09391_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[17] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[18] ),
    .C(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__mux4_1 _09392_ (.A0(_03697_),
    .A1(_03698_),
    .A2(_03786_),
    .A3(_03787_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ),
    .X(_03840_));
 sky130_fd_sc_hd__inv_2 _09393_ (.A(net3677),
    .Y(_03841_));
 sky130_fd_sc_hd__o31a_1 _09394_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[17] ),
    .A2(_03833_),
    .A3(_03840_),
    .B1(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__mux4_1 _09395_ (.A0(_03484_),
    .A1(_03486_),
    .A2(_03488_),
    .A3(_03490_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ),
    .X(_03843_));
 sky130_fd_sc_hd__inv_2 _09396_ (.A(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__mux4_1 _09397_ (.A0(_03503_),
    .A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ),
    .X(_03845_));
 sky130_fd_sc_hd__mux4_1 _09398_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ),
    .X(_03846_));
 sky130_fd_sc_hd__and3b_1 _09399_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[17] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[18] ),
    .C(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__a31oi_1 _09400_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[17] ),
    .A2(_03833_),
    .A3(_03845_),
    .B1(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__o311a_1 _09401_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[17] ),
    .A2(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[18] ),
    .A3(_03844_),
    .B1(_03848_),
    .C1(net3677),
    .X(_03849_));
 sky130_fd_sc_hd__a31oi_1 _09402_ (.A1(_03837_),
    .A2(_03839_),
    .A3(net3678),
    .B1(_03849_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[3] ));
 sky130_fd_sc_hd__mux4_1 _09403_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ),
    .X(_03850_));
 sky130_fd_sc_hd__mux4_1 _09404_ (.A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ),
    .X(_03851_));
 sky130_fd_sc_hd__o21ai_1 _09405_ (.A1(_00359_),
    .A2(_03851_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[12] ),
    .Y(_03852_));
 sky130_fd_sc_hd__a21oi_1 _09406_ (.A1(_00359_),
    .A2(_03850_),
    .B1(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hd__nor2_1 _09407_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[12] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[13] ),
    .Y(_03854_));
 sky130_fd_sc_hd__mux4_1 _09408_ (.A0(_03780_),
    .A1(_03781_),
    .A2(_03782_),
    .A3(_03783_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ),
    .S1(_00351_),
    .X(_03855_));
 sky130_fd_sc_hd__and2_1 _09409_ (.A(_03854_),
    .B(_03855_),
    .X(_03856_));
 sky130_fd_sc_hd__mux4_1 _09410_ (.A0(_03530_),
    .A1(_03531_),
    .A2(_03786_),
    .A3(_03787_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ),
    .X(_03857_));
 sky130_fd_sc_hd__nor3_1 _09411_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[12] ),
    .B(_00359_),
    .C(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__mux4_1 _09412_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ),
    .X(_03859_));
 sky130_fd_sc_hd__mux4_1 _09413_ (.A0(_03494_),
    .A1(_03496_),
    .A2(_03498_),
    .A3(_03500_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ),
    .X(_03860_));
 sky130_fd_sc_hd__and3_1 _09414_ (.A(_00355_),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[13] ),
    .C(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__mux4_1 _09415_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ),
    .X(_03862_));
 sky130_fd_sc_hd__a31o_1 _09416_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[12] ),
    .A2(_00359_),
    .A3(_03862_),
    .B1(_00361_),
    .X(_03863_));
 sky130_fd_sc_hd__a211o_1 _09417_ (.A1(_03854_),
    .A2(_03859_),
    .B1(_03861_),
    .C1(_03863_),
    .X(_03864_));
 sky130_fd_sc_hd__o41a_1 _09418_ (.A1(net3168),
    .A2(_03853_),
    .A3(_03856_),
    .A4(net3246),
    .B1(_03864_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[2] ));
 sky130_fd_sc_hd__clkbuf_4 _09419_ (.A(_00171_),
    .X(_03865_));
 sky130_fd_sc_hd__nand3b_2 _09420_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .C(_01415_),
    .Y(_03866_));
 sky130_fd_sc_hd__or3_1 _09421_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_03867_));
 sky130_fd_sc_hd__or2_1 _09422_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__clkbuf_2 _09423_ (.A(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__o21a_2 _09424_ (.A1(_03866_),
    .A2(_03869_),
    .B1(_03013_),
    .X(_03870_));
 sky130_fd_sc_hd__mux2_1 _09425_ (.A0(_03865_),
    .A1(net3603),
    .S(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__clkbuf_1 _09426_ (.A(_03871_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__clkbuf_4 _09427_ (.A(_00184_),
    .X(_03872_));
 sky130_fd_sc_hd__mux2_1 _09428_ (.A0(_03872_),
    .A1(net3467),
    .S(_03870_),
    .X(_03873_));
 sky130_fd_sc_hd__clkbuf_1 _09429_ (.A(_03873_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__clkbuf_4 _09430_ (.A(_00551_),
    .X(_03874_));
 sky130_fd_sc_hd__mux2_1 _09431_ (.A0(_03874_),
    .A1(net3436),
    .S(_03870_),
    .X(_03875_));
 sky130_fd_sc_hd__clkbuf_1 _09432_ (.A(_03875_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _09433_ (.A0(_03622_),
    .A1(net3444),
    .S(_03870_),
    .X(_03876_));
 sky130_fd_sc_hd__clkbuf_1 _09434_ (.A(_03876_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__buf_2 _09435_ (.A(net4048),
    .X(_03877_));
 sky130_fd_sc_hd__clkbuf_2 _09436_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ),
    .X(_03878_));
 sky130_fd_sc_hd__inv_2 _09437_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .Y(_03879_));
 sky130_fd_sc_hd__or4_1 _09438_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03878_),
    .C(_03879_),
    .D(_03866_),
    .X(_03880_));
 sky130_fd_sc_hd__o21a_2 _09439_ (.A1(_03877_),
    .A2(_03880_),
    .B1(_01489_),
    .X(_03881_));
 sky130_fd_sc_hd__mux2_1 _09440_ (.A0(_03865_),
    .A1(net3531),
    .S(_03881_),
    .X(_03882_));
 sky130_fd_sc_hd__clkbuf_1 _09441_ (.A(_03882_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _09442_ (.A0(_03872_),
    .A1(net3547),
    .S(_03881_),
    .X(_03883_));
 sky130_fd_sc_hd__clkbuf_1 _09443_ (.A(_03883_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _09444_ (.A0(_03874_),
    .A1(net3479),
    .S(_03881_),
    .X(_03884_));
 sky130_fd_sc_hd__clkbuf_1 _09445_ (.A(_03884_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _09446_ (.A0(_03622_),
    .A1(net3342),
    .S(_03881_),
    .X(_03885_));
 sky130_fd_sc_hd__clkbuf_1 _09447_ (.A(_03885_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__mux4_1 _09448_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ),
    .X(_03886_));
 sky130_fd_sc_hd__mux4_1 _09449_ (.A0(_03816_),
    .A1(_03817_),
    .A2(_03818_),
    .A3(_03819_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ),
    .X(_03887_));
 sky130_fd_sc_hd__nor2_1 _09450_ (.A(_00344_),
    .B(_03887_),
    .Y(_03888_));
 sky130_fd_sc_hd__a211o_1 _09451_ (.A1(_00344_),
    .A2(_03886_),
    .B1(_03888_),
    .C1(_00342_),
    .X(_03889_));
 sky130_fd_sc_hd__mux4_1 _09452_ (.A0(_00784_),
    .A1(_01143_),
    .A2(_01227_),
    .A3(_01056_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ),
    .S1(_00336_),
    .X(_03890_));
 sky130_fd_sc_hd__or3_1 _09453_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[7] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[8] ),
    .C(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__mux4_1 _09454_ (.A0(_03697_),
    .A1(_03698_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ),
    .X(_03892_));
 sky130_fd_sc_hd__o31a_1 _09455_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[7] ),
    .A2(_00344_),
    .A3(_03892_),
    .B1(_00349_),
    .X(_03893_));
 sky130_fd_sc_hd__mux4_1 _09456_ (.A0(_03484_),
    .A1(_03486_),
    .A2(_03488_),
    .A3(_03490_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ),
    .X(_03894_));
 sky130_fd_sc_hd__mux4_1 _09457_ (.A0(_03806_),
    .A1(_03807_),
    .A2(_03808_),
    .A3(_03809_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ),
    .X(_03895_));
 sky130_fd_sc_hd__mux4_1 _09458_ (.A0(_03493_),
    .A1(_03495_),
    .A2(_03497_),
    .A3(_03499_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ),
    .X(_03896_));
 sky130_fd_sc_hd__and3_1 _09459_ (.A(_00342_),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[8] ),
    .C(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__a31o_1 _09460_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[7] ),
    .A2(_00344_),
    .A3(_03895_),
    .B1(_03897_),
    .X(_03898_));
 sky130_fd_sc_hd__a311oi_1 _09461_ (.A1(_00342_),
    .A2(_00344_),
    .A3(_03894_),
    .B1(_03898_),
    .C1(_00349_),
    .Y(_03899_));
 sky130_fd_sc_hd__a31oi_1 _09462_ (.A1(_03889_),
    .A2(_03891_),
    .A3(_03893_),
    .B1(net3619),
    .Y(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[1] ));
 sky130_fd_sc_hd__inv_2 _09463_ (.A(_03877_),
    .Y(_03900_));
 sky130_fd_sc_hd__or3_2 _09464_ (.A(_03878_),
    .B(_03900_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_03901_));
 sky130_fd_sc_hd__and3b_1 _09465_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .C(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ),
    .X(_03902_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09466_ (.A(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__nand2_1 _09467_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03867_),
    .Y(_03904_));
 sky130_fd_sc_hd__and2_1 _09468_ (.A(_03869_),
    .B(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__nand2_1 _09469_ (.A(_03903_),
    .B(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__nand2_1 _09470_ (.A(_02003_),
    .B(_03869_),
    .Y(_03907_));
 sky130_fd_sc_hd__or3_1 _09471_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03866_),
    .C(_03901_),
    .X(_03908_));
 sky130_fd_sc_hd__nand2_1 _09472_ (.A(net3785),
    .B(_03908_),
    .Y(_03909_));
 sky130_fd_sc_hd__o31a_1 _09473_ (.A1(_03901_),
    .A2(_03906_),
    .A3(_03907_),
    .B1(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__o21ai_1 _09474_ (.A1(_03408_),
    .A2(_03910_),
    .B1(_02978_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_2 _09475_ (.A(_01446_),
    .B(_03869_),
    .Y(_03911_));
 sky130_fd_sc_hd__nand2_1 _09476_ (.A(net3351),
    .B(_03908_),
    .Y(_03912_));
 sky130_fd_sc_hd__o31a_1 _09477_ (.A1(_03901_),
    .A2(_03906_),
    .A3(_03911_),
    .B1(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__o21ai_1 _09478_ (.A1(_03408_),
    .A2(_03913_),
    .B1(_03379_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__clkbuf_4 _09479_ (.A(_01764_),
    .X(_03914_));
 sky130_fd_sc_hd__nand2_1 _09480_ (.A(_02573_),
    .B(_03869_),
    .Y(_03915_));
 sky130_fd_sc_hd__nand2_1 _09481_ (.A(net3723),
    .B(_03908_),
    .Y(_03916_));
 sky130_fd_sc_hd__o31a_1 _09482_ (.A1(_03901_),
    .A2(_03906_),
    .A3(_03915_),
    .B1(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__o21ai_1 _09483_ (.A1(_03914_),
    .A2(_03917_),
    .B1(_00251_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__nand2_1 _09484_ (.A(_00264_),
    .B(_03869_),
    .Y(_03918_));
 sky130_fd_sc_hd__nand2_1 _09485_ (.A(net3812),
    .B(_03908_),
    .Y(_03919_));
 sky130_fd_sc_hd__o31a_1 _09486_ (.A1(_03901_),
    .A2(_03906_),
    .A3(_03918_),
    .B1(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__o21ai_1 _09487_ (.A1(_03914_),
    .A2(_03920_),
    .B1(_03322_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _09488_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03866_),
    .Y(_03921_));
 sky130_fd_sc_hd__and3b_1 _09489_ (.A_N(_03878_),
    .B(_03877_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(_03922_));
 sky130_fd_sc_hd__a21oi_4 _09490_ (.A1(_03921_),
    .A2(_03922_),
    .B1(_02686_),
    .Y(_03923_));
 sky130_fd_sc_hd__mux2_1 _09491_ (.A0(_03865_),
    .A1(net3487),
    .S(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__clkbuf_1 _09492_ (.A(_03924_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _09493_ (.A0(_03872_),
    .A1(net3350),
    .S(_03923_),
    .X(_03925_));
 sky130_fd_sc_hd__clkbuf_1 _09494_ (.A(_03925_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _09495_ (.A0(_03874_),
    .A1(net3460),
    .S(_03923_),
    .X(_03926_));
 sky130_fd_sc_hd__clkbuf_1 _09496_ (.A(_03926_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _09497_ (.A0(_03622_),
    .A1(net3483),
    .S(_03923_),
    .X(_03927_));
 sky130_fd_sc_hd__clkbuf_1 _09498_ (.A(_03927_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4_1 _09499_ (.A(_03878_),
    .B(_03900_),
    .C(_03879_),
    .D(_03921_),
    .X(_03928_));
 sky130_fd_sc_hd__clkbuf_2 _09500_ (.A(_03928_),
    .X(_03929_));
 sky130_fd_sc_hd__nand2_1 _09501_ (.A(_03907_),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__or2_1 _09502_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .B(_03929_),
    .X(_03931_));
 sky130_fd_sc_hd__a31o_1 _09503_ (.A1(_03666_),
    .A2(_03930_),
    .A3(_03931_),
    .B1(_03316_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _09504_ (.A(_03911_),
    .B(_03929_),
    .Y(_03932_));
 sky130_fd_sc_hd__or2_1 _09505_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .B(_03929_),
    .X(_03933_));
 sky130_fd_sc_hd__a31o_1 _09506_ (.A1(_03666_),
    .A2(_03932_),
    .A3(_03933_),
    .B1(_01772_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _09507_ (.A(_03915_),
    .B(_03929_),
    .Y(_03934_));
 sky130_fd_sc_hd__or2_1 _09508_ (.A(net4081),
    .B(_03929_),
    .X(_03935_));
 sky130_fd_sc_hd__a31o_1 _09509_ (.A1(_03666_),
    .A2(_03934_),
    .A3(_03935_),
    .B1(_01851_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _09510_ (.A(net3972),
    .B(_03929_),
    .Y(_03936_));
 sky130_fd_sc_hd__a211o_1 _09511_ (.A1(_03918_),
    .A2(_03929_),
    .B1(_03936_),
    .C1(_00228_),
    .X(_03937_));
 sky130_fd_sc_hd__nand2_1 _09512_ (.A(_03166_),
    .B(_03937_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _09513_ (.A1(_03878_),
    .A2(_03900_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .A4(_03921_),
    .B1(_00249_),
    .X(_03938_));
 sky130_fd_sc_hd__mux2_1 _09514_ (.A0(net4013),
    .A1(_03169_),
    .S(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__clkbuf_1 _09515_ (.A(_03939_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _09516_ (.A0(net4187),
    .A1(_03172_),
    .S(_03938_),
    .X(_03940_));
 sky130_fd_sc_hd__clkbuf_1 _09517_ (.A(_03940_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__inv_2 _09518_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[3] ),
    .Y(_03941_));
 sky130_fd_sc_hd__mux4_1 _09519_ (.A0(_03511_),
    .A1(_03512_),
    .A2(_03513_),
    .A3(_03514_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[1] ),
    .X(_03942_));
 sky130_fd_sc_hd__mux4_1 _09520_ (.A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[1] ),
    .X(_03943_));
 sky130_fd_sc_hd__o21ai_1 _09521_ (.A1(_03941_),
    .A2(_03943_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[2] ),
    .Y(_03944_));
 sky130_fd_sc_hd__a21oi_1 _09522_ (.A1(_03941_),
    .A2(_03942_),
    .B1(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__mux4_1 _09523_ (.A0(_03530_),
    .A1(_03531_),
    .A2(_03532_),
    .A3(_03533_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[1] ),
    .X(_03946_));
 sky130_fd_sc_hd__nor3_1 _09524_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[2] ),
    .B(_03941_),
    .C(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__mux4_1 _09525_ (.A0(_03758_),
    .A1(_03759_),
    .A2(_03760_),
    .A3(_03761_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[1] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[0] ),
    .X(_03948_));
 sky130_fd_sc_hd__o31ai_1 _09526_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[2] ),
    .A2(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[3] ),
    .A3(_03948_),
    .B1(_00332_),
    .Y(_03949_));
 sky130_fd_sc_hd__nor2_1 _09527_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[2] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[3] ),
    .Y(_03950_));
 sky130_fd_sc_hd__mux4_1 _09528_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[1] ),
    .X(_03951_));
 sky130_fd_sc_hd__mux4_1 _09529_ (.A0(_03494_),
    .A1(_03496_),
    .A2(_03498_),
    .A3(_03500_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[1] ),
    .X(_03952_));
 sky130_fd_sc_hd__and3b_1 _09530_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[2] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[3] ),
    .C(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__mux4_1 _09531_ (.A0(_03503_),
    .A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[1] ),
    .X(_03954_));
 sky130_fd_sc_hd__a31o_1 _09532_ (.A1(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[2] ),
    .A2(_03941_),
    .A3(_03954_),
    .B1(_00332_),
    .X(_03955_));
 sky130_fd_sc_hd__a211o_1 _09533_ (.A1(_03950_),
    .A2(_03951_),
    .B1(_03953_),
    .C1(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__o31a_1 _09534_ (.A1(_03945_),
    .A2(_03947_),
    .A3(_03949_),
    .B1(_03956_),
    .X(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[0] ));
 sky130_fd_sc_hd__mux2_1 _09535_ (.A0(net4023),
    .A1(_03174_),
    .S(_03938_),
    .X(_03957_));
 sky130_fd_sc_hd__clkbuf_1 _09536_ (.A(_03957_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _09537_ (.A0(net3760),
    .A1(_00527_),
    .S(_03938_),
    .X(_03958_));
 sky130_fd_sc_hd__clkbuf_1 _09538_ (.A(_03958_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_1 _09539_ (.A(_03878_),
    .B(_03877_),
    .C(_03879_),
    .D(_03921_),
    .X(_03959_));
 sky130_fd_sc_hd__or2_1 _09540_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .B(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__nand2_1 _09541_ (.A(_03907_),
    .B(_03959_),
    .Y(_03961_));
 sky130_fd_sc_hd__a31o_1 _09542_ (.A1(_03666_),
    .A2(_03960_),
    .A3(_03961_),
    .B1(_03316_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _09543_ (.A0(_00715_),
    .A1(_03911_),
    .S(_03959_),
    .X(_03962_));
 sky130_fd_sc_hd__o21ai_1 _09544_ (.A1(_03914_),
    .A2(_03962_),
    .B1(_03379_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _09545_ (.A0(_00722_),
    .A1(_03915_),
    .S(_03959_),
    .X(_03963_));
 sky130_fd_sc_hd__o21ai_1 _09546_ (.A1(_03914_),
    .A2(_03963_),
    .B1(_00251_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _09547_ (.A0(_00718_),
    .A1(_03918_),
    .S(_03959_),
    .X(_03964_));
 sky130_fd_sc_hd__o21ai_1 _09548_ (.A1(_03914_),
    .A2(_03964_),
    .B1(_03322_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _09549_ (.A1(_03878_),
    .A2(_03877_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .A4(_03921_),
    .B1(_00249_),
    .X(_03965_));
 sky130_fd_sc_hd__mux2_1 _09550_ (.A0(net4087),
    .A1(_03169_),
    .S(_03965_),
    .X(_03966_));
 sky130_fd_sc_hd__clkbuf_1 _09551_ (.A(_03966_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _09552_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .A1(_03172_),
    .S(_03965_),
    .X(_03967_));
 sky130_fd_sc_hd__clkbuf_1 _09553_ (.A(_03967_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _09554_ (.A0(net3822),
    .A1(_03174_),
    .S(_03965_),
    .X(_03968_));
 sky130_fd_sc_hd__clkbuf_1 _09555_ (.A(_03968_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _09556_ (.A0(net4181),
    .A1(_00527_),
    .S(_03965_),
    .X(_03969_));
 sky130_fd_sc_hd__clkbuf_1 _09557_ (.A(_03969_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _09558_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .Y(_03970_));
 sky130_fd_sc_hd__o31a_2 _09559_ (.A1(_03970_),
    .A2(_03866_),
    .A3(_03867_),
    .B1(_02847_),
    .X(_03971_));
 sky130_fd_sc_hd__mux2_1 _09560_ (.A0(_03865_),
    .A1(net3855),
    .S(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__clkbuf_1 _09561_ (.A(_03972_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _09562_ (.A0(_03872_),
    .A1(net3403),
    .S(_03971_),
    .X(_03973_));
 sky130_fd_sc_hd__clkbuf_1 _09563_ (.A(_03973_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _09564_ (.A0(_03874_),
    .A1(net3596),
    .S(_03971_),
    .X(_03974_));
 sky130_fd_sc_hd__clkbuf_1 _09565_ (.A(_03974_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _09566_ (.A0(_03622_),
    .A1(net3840),
    .S(_03971_),
    .X(_03975_));
 sky130_fd_sc_hd__clkbuf_1 _09567_ (.A(_03975_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _09568_ (.A(_03866_),
    .B(_03905_),
    .X(_03976_));
 sky130_fd_sc_hd__o41a_2 _09569_ (.A1(_03878_),
    .A2(_03877_),
    .A3(_03879_),
    .A4(_03976_),
    .B1(_00407_),
    .X(_03977_));
 sky130_fd_sc_hd__mux2_1 _09570_ (.A0(_03865_),
    .A1(net3660),
    .S(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__clkbuf_1 _09571_ (.A(_03978_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _09572_ (.A0(_03872_),
    .A1(net3707),
    .S(_03977_),
    .X(_03979_));
 sky130_fd_sc_hd__clkbuf_1 _09573_ (.A(_03979_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _09574_ (.A0(_03874_),
    .A1(net3708),
    .S(_03977_),
    .X(_03980_));
 sky130_fd_sc_hd__clkbuf_1 _09575_ (.A(_03980_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _09576_ (.A0(_03622_),
    .A1(net3691),
    .S(_03977_),
    .X(_03981_));
 sky130_fd_sc_hd__clkbuf_1 _09577_ (.A(_03981_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__clkbuf_4 _09578_ (.A(_00195_),
    .X(_03982_));
 sky130_fd_sc_hd__nor2_2 _09579_ (.A(_03901_),
    .B(_03976_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _09580_ (.A(_03907_),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__or2_1 _09581_ (.A(net4109),
    .B(_03983_),
    .X(_03985_));
 sky130_fd_sc_hd__a31o_1 _09582_ (.A1(_03982_),
    .A2(_03984_),
    .A3(_03985_),
    .B1(_03316_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__mux2_1 _09583_ (.A0(_03211_),
    .A1(_03911_),
    .S(_03983_),
    .X(_03986_));
 sky130_fd_sc_hd__o21ai_1 _09584_ (.A1(_03914_),
    .A2(_03986_),
    .B1(_03379_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__mux2_1 _09585_ (.A0(_03214_),
    .A1(_03915_),
    .S(_03983_),
    .X(_03987_));
 sky130_fd_sc_hd__o21ai_1 _09586_ (.A1(_03914_),
    .A2(_03987_),
    .B1(_00251_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__nor2_1 _09587_ (.A(net3400),
    .B(_03983_),
    .Y(_03988_));
 sky130_fd_sc_hd__a211o_1 _09588_ (.A1(_03918_),
    .A2(_03983_),
    .B1(_03988_),
    .C1(_00228_),
    .X(_03989_));
 sky130_fd_sc_hd__nand2_1 _09589_ (.A(_03166_),
    .B(_03989_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3_2 _09590_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(_03903_),
    .C(_03922_),
    .X(_03990_));
 sky130_fd_sc_hd__nor2_1 _09591_ (.A(_01971_),
    .B(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__a221o_1 _09592_ (.A1(_00288_),
    .A2(_03990_),
    .B1(_03991_),
    .B2(net3158),
    .C1(_00209_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _09593_ (.A1(_00293_),
    .A2(_03990_),
    .B1(_03991_),
    .B2(net3133),
    .C1(_02872_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _09594_ (.A1(_00295_),
    .A2(_03990_),
    .B1(_03991_),
    .B2(net3250),
    .C1(_00221_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__and2_1 _09595_ (.A(_01578_),
    .B(_00781_),
    .X(_03992_));
 sky130_fd_sc_hd__buf_4 _09596_ (.A(_01862_),
    .X(_03993_));
 sky130_fd_sc_hd__mux2_1 _09597_ (.A0(_03751_),
    .A1(_03992_),
    .S(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__clkbuf_1 _09598_ (.A(_03994_),
    .X(_00001_));
 sky130_fd_sc_hd__mux4_1 _09599_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[36] ),
    .X(_03995_));
 sky130_fd_sc_hd__mux4_1 _09600_ (.A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[36] ),
    .X(_03996_));
 sky130_fd_sc_hd__o21a_1 _09601_ (.A1(_00536_),
    .A2(_03996_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[37] ),
    .X(_03997_));
 sky130_fd_sc_hd__o21ai_1 _09602_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[38] ),
    .A2(_03995_),
    .B1(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hd__mux4_1 _09603_ (.A0(_03759_),
    .A1(_03758_),
    .A2(_03761_),
    .A3(_03760_),
    .S0(_00532_),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ),
    .X(_03999_));
 sky130_fd_sc_hd__o31a_1 _09604_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[37] ),
    .A2(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[38] ),
    .A3(_03999_),
    .B1(_00538_),
    .X(_04000_));
 sky130_fd_sc_hd__mux4_1 _09605_ (.A0(_03697_),
    .A1(_03698_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[36] ),
    .X(_04001_));
 sky130_fd_sc_hd__or3_1 _09606_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[37] ),
    .B(_00536_),
    .C(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__mux4_1 _09607_ (.A0(_03806_),
    .A1(_03807_),
    .A2(_03808_),
    .A3(_03809_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[36] ),
    .X(_04003_));
 sky130_fd_sc_hd__a31o_1 _09608_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[37] ),
    .A2(_00536_),
    .A3(_04003_),
    .B1(_00538_),
    .X(_04004_));
 sky130_fd_sc_hd__mux4_1 _09609_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[36] ),
    .X(_04005_));
 sky130_fd_sc_hd__or3b_1 _09610_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[37] ),
    .B(_00536_),
    .C_N(_04005_),
    .X(_04006_));
 sky130_fd_sc_hd__mux4_1 _09611_ (.A0(net21),
    .A1(net22),
    .A2(net23),
    .A3(net24),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[36] ),
    .X(_04007_));
 sky130_fd_sc_hd__or3b_1 _09612_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[37] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[38] ),
    .C_N(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__and3b_1 _09613_ (.A_N(_04004_),
    .B(_04006_),
    .C(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__a31oi_1 _09614_ (.A1(_03998_),
    .A2(net3505),
    .A3(_04002_),
    .B1(_04009_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[7] ));
 sky130_fd_sc_hd__mux4_1 _09615_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[31] ),
    .X(_04010_));
 sky130_fd_sc_hd__inv_2 _09616_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ),
    .Y(_04011_));
 sky130_fd_sc_hd__mux4_1 _09617_ (.A0(_03816_),
    .A1(_03817_),
    .A2(_03818_),
    .A3(_03819_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[31] ),
    .X(_04012_));
 sky130_fd_sc_hd__or2_1 _09618_ (.A(_04011_),
    .B(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__o211a_1 _09619_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ),
    .A2(_04010_),
    .B1(_04013_),
    .C1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ),
    .X(_04014_));
 sky130_fd_sc_hd__mux4_1 _09620_ (.A0(_03530_),
    .A1(_03531_),
    .A2(_03532_),
    .A3(_03533_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[31] ),
    .X(_04015_));
 sky130_fd_sc_hd__nor3_1 _09621_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ),
    .B(_04011_),
    .C(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__nor2_1 _09622_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ),
    .Y(_04017_));
 sky130_fd_sc_hd__mux4_1 _09623_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[31] ),
    .S1(_00518_),
    .X(_04018_));
 sky130_fd_sc_hd__a21o_1 _09624_ (.A1(_04017_),
    .A2(_04018_),
    .B1(net3999),
    .X(_04019_));
 sky130_fd_sc_hd__mux4_1 _09625_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[31] ),
    .X(_04020_));
 sky130_fd_sc_hd__mux4_1 _09626_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[31] ),
    .X(_04021_));
 sky130_fd_sc_hd__mux4_1 _09627_ (.A0(_03493_),
    .A1(_03495_),
    .A2(_03497_),
    .A3(_03499_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[31] ),
    .X(_04022_));
 sky130_fd_sc_hd__and3b_1 _09628_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ),
    .C(_04022_),
    .X(_04023_));
 sky130_fd_sc_hd__a31o_1 _09629_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ),
    .A2(_04011_),
    .A3(_04021_),
    .B1(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__inv_2 _09630_ (.A(net3999),
    .Y(_04025_));
 sky130_fd_sc_hd__a211o_1 _09631_ (.A1(_04017_),
    .A2(_04020_),
    .B1(_04024_),
    .C1(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__o31a_1 _09632_ (.A1(_04014_),
    .A2(_04016_),
    .A3(_04019_),
    .B1(_04026_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[6] ));
 sky130_fd_sc_hd__mux4_1 _09633_ (.A0(_02226_),
    .A1(_02320_),
    .A2(_02408_),
    .A3(_02491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[26] ),
    .X(_04027_));
 sky130_fd_sc_hd__mux4_1 _09634_ (.A0(_03816_),
    .A1(_03817_),
    .A2(_03818_),
    .A3(_03819_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[26] ),
    .X(_04028_));
 sky130_fd_sc_hd__or2_1 _09635_ (.A(_00513_),
    .B(_04028_),
    .X(_04029_));
 sky130_fd_sc_hd__o211a_1 _09636_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[28] ),
    .A2(_04027_),
    .B1(_04029_),
    .C1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[27] ),
    .X(_04030_));
 sky130_fd_sc_hd__nor2_1 _09637_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[27] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[28] ),
    .Y(_04031_));
 sky130_fd_sc_hd__mux4_1 _09638_ (.A0(_03780_),
    .A1(_03781_),
    .A2(_03782_),
    .A3(_03783_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[26] ),
    .S1(_00506_),
    .X(_04032_));
 sky130_fd_sc_hd__and2_1 _09639_ (.A(_04031_),
    .B(_04032_),
    .X(_04033_));
 sky130_fd_sc_hd__mux4_1 _09640_ (.A0(_03530_),
    .A1(_03531_),
    .A2(_03786_),
    .A3(_03787_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[26] ),
    .X(_04034_));
 sky130_fd_sc_hd__nor3_1 _09641_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[27] ),
    .B(_00513_),
    .C(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__mux4_1 _09642_ (.A0(_03485_),
    .A1(_03487_),
    .A2(_03489_),
    .A3(_03491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[26] ),
    .X(_04036_));
 sky130_fd_sc_hd__mux4_1 _09643_ (.A0(_03494_),
    .A1(_03496_),
    .A2(_03498_),
    .A3(_03500_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[26] ),
    .X(_04037_));
 sky130_fd_sc_hd__and3_1 _09644_ (.A(_00511_),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[28] ),
    .C(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__mux4_1 _09645_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[26] ),
    .X(_04039_));
 sky130_fd_sc_hd__a31o_1 _09646_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[27] ),
    .A2(_00513_),
    .A3(_04039_),
    .B1(_00516_),
    .X(_04040_));
 sky130_fd_sc_hd__a211o_1 _09647_ (.A1(_04031_),
    .A2(_04036_),
    .B1(_04038_),
    .C1(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__o41a_1 _09648_ (.A1(net3309),
    .A2(_04030_),
    .A3(_04033_),
    .A4(_04035_),
    .B1(_04041_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[5] ));
 sky130_fd_sc_hd__mux4_1 _09649_ (.A0(_02226_),
    .A1(_02320_),
    .A2(_02408_),
    .A3(_02491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[21] ),
    .X(_04042_));
 sky130_fd_sc_hd__mux4_1 _09650_ (.A0(_03816_),
    .A1(_03817_),
    .A2(_03818_),
    .A3(_03819_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[21] ),
    .X(_04043_));
 sky130_fd_sc_hd__or2_1 _09651_ (.A(_00500_),
    .B(_04043_),
    .X(_04044_));
 sky130_fd_sc_hd__o211a_1 _09652_ (.A1(net4224),
    .A2(_04042_),
    .B1(_04044_),
    .C1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[22] ),
    .X(_04045_));
 sky130_fd_sc_hd__nor2_1 _09653_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[22] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[23] ),
    .Y(_04046_));
 sky130_fd_sc_hd__mux4_1 _09654_ (.A0(_03780_),
    .A1(_03781_),
    .A2(_03782_),
    .A3(_03783_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[21] ),
    .S1(_00492_),
    .X(_04047_));
 sky130_fd_sc_hd__and2_1 _09655_ (.A(_04046_),
    .B(_04047_),
    .X(_04048_));
 sky130_fd_sc_hd__mux4_1 _09656_ (.A0(_03530_),
    .A1(_03531_),
    .A2(_03786_),
    .A3(_03787_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[21] ),
    .X(_04049_));
 sky130_fd_sc_hd__nor3_1 _09657_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[22] ),
    .B(_00500_),
    .C(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__mux4_1 _09658_ (.A0(_03485_),
    .A1(_03487_),
    .A2(_03489_),
    .A3(_03491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[21] ),
    .X(_04051_));
 sky130_fd_sc_hd__mux4_1 _09659_ (.A0(_03494_),
    .A1(_03496_),
    .A2(_03498_),
    .A3(_03500_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[21] ),
    .X(_04052_));
 sky130_fd_sc_hd__and3_1 _09660_ (.A(_00498_),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[23] ),
    .C(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__mux4_1 _09661_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[21] ),
    .X(_04054_));
 sky130_fd_sc_hd__a31o_1 _09662_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[22] ),
    .A2(_00500_),
    .A3(_04054_),
    .B1(_00502_),
    .X(_04055_));
 sky130_fd_sc_hd__a211o_1 _09663_ (.A1(_04046_),
    .A2(_04051_),
    .B1(_04053_),
    .C1(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__o41a_1 _09664_ (.A1(net3256),
    .A2(net4225),
    .A3(_04048_),
    .A4(_04050_),
    .B1(_04056_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[4] ));
 sky130_fd_sc_hd__mux4_1 _09665_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[16] ),
    .X(_04057_));
 sky130_fd_sc_hd__inv_2 _09666_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[18] ),
    .Y(_04058_));
 sky130_fd_sc_hd__mux4_1 _09667_ (.A0(_03816_),
    .A1(_03817_),
    .A2(_03818_),
    .A3(_03819_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[16] ),
    .X(_04059_));
 sky130_fd_sc_hd__or2_1 _09668_ (.A(_04058_),
    .B(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__o211a_1 _09669_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[18] ),
    .A2(_04057_),
    .B1(_04060_),
    .C1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[17] ),
    .X(_04061_));
 sky130_fd_sc_hd__mux4_1 _09670_ (.A0(_03530_),
    .A1(_03531_),
    .A2(_03532_),
    .A3(_03533_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[16] ),
    .X(_04062_));
 sky130_fd_sc_hd__nor3_1 _09671_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[17] ),
    .B(_04058_),
    .C(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__nor2_1 _09672_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[17] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[18] ),
    .Y(_04064_));
 sky130_fd_sc_hd__mux4_1 _09673_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[16] ),
    .S1(_00480_),
    .X(_04065_));
 sky130_fd_sc_hd__a21o_1 _09674_ (.A1(_04064_),
    .A2(_04065_),
    .B1(net3433),
    .X(_04066_));
 sky130_fd_sc_hd__mux4_1 _09675_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[16] ),
    .X(_04067_));
 sky130_fd_sc_hd__mux4_1 _09676_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[16] ),
    .X(_04068_));
 sky130_fd_sc_hd__mux4_1 _09677_ (.A0(_03493_),
    .A1(_03495_),
    .A2(_03497_),
    .A3(_03499_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[16] ),
    .X(_04069_));
 sky130_fd_sc_hd__and3b_1 _09678_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[17] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[18] ),
    .C(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__a31o_1 _09679_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[17] ),
    .A2(_04058_),
    .A3(_04068_),
    .B1(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__inv_2 _09680_ (.A(net3433),
    .Y(_04072_));
 sky130_fd_sc_hd__a211o_1 _09681_ (.A1(_04064_),
    .A2(_04067_),
    .B1(_04071_),
    .C1(_04072_),
    .X(_04073_));
 sky130_fd_sc_hd__o31a_1 _09682_ (.A1(_04061_),
    .A2(_04063_),
    .A3(_04066_),
    .B1(_04073_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[3] ));
 sky130_fd_sc_hd__mux4_1 _09683_ (.A0(_02226_),
    .A1(_02320_),
    .A2(_02408_),
    .A3(_02491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ),
    .X(_04074_));
 sky130_fd_sc_hd__mux4_1 _09684_ (.A0(_03816_),
    .A1(_03817_),
    .A2(_03818_),
    .A3(_03819_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ),
    .X(_04075_));
 sky130_fd_sc_hd__or2_1 _09685_ (.A(_00475_),
    .B(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__o211a_1 _09686_ (.A1(net4231),
    .A2(_04074_),
    .B1(_04076_),
    .C1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[12] ),
    .X(_04077_));
 sky130_fd_sc_hd__nor2_1 _09687_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[12] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[13] ),
    .Y(_04078_));
 sky130_fd_sc_hd__mux4_1 _09688_ (.A0(_03780_),
    .A1(_03781_),
    .A2(_03782_),
    .A3(_03783_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ),
    .S1(_00467_),
    .X(_04079_));
 sky130_fd_sc_hd__and2_1 _09689_ (.A(_04078_),
    .B(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__mux4_1 _09690_ (.A0(_03697_),
    .A1(_03531_),
    .A2(_03786_),
    .A3(_03787_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ),
    .X(_04081_));
 sky130_fd_sc_hd__nor3_1 _09691_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[12] ),
    .B(_00475_),
    .C(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__mux4_1 _09692_ (.A0(_03485_),
    .A1(_03487_),
    .A2(_03489_),
    .A3(_03491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ),
    .X(_04083_));
 sky130_fd_sc_hd__mux4_1 _09693_ (.A0(_03494_),
    .A1(_03496_),
    .A2(_03498_),
    .A3(_03500_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ),
    .X(_04084_));
 sky130_fd_sc_hd__and3_1 _09694_ (.A(_00471_),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[13] ),
    .C(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__mux4_1 _09695_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ),
    .X(_04086_));
 sky130_fd_sc_hd__a31o_1 _09696_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[12] ),
    .A2(_00475_),
    .A3(_04086_),
    .B1(_00477_),
    .X(_04087_));
 sky130_fd_sc_hd__a211o_1 _09697_ (.A1(_04078_),
    .A2(_04083_),
    .B1(_04085_),
    .C1(_04087_),
    .X(_04088_));
 sky130_fd_sc_hd__o41a_1 _09698_ (.A1(net3395),
    .A2(_04077_),
    .A3(_04080_),
    .A4(_04082_),
    .B1(_04088_),
    .X(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[2] ));
 sky130_fd_sc_hd__mux4_1 _09699_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ),
    .X(_04089_));
 sky130_fd_sc_hd__mux4_1 _09700_ (.A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ),
    .X(_04090_));
 sky130_fd_sc_hd__o21a_1 _09701_ (.A1(_00458_),
    .A2(_04090_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[7] ),
    .X(_04091_));
 sky130_fd_sc_hd__o21ai_1 _09702_ (.A1(net3422),
    .A2(_04089_),
    .B1(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__mux4_1 _09703_ (.A0(_03760_),
    .A1(_03761_),
    .A2(_03758_),
    .A3(_03759_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ),
    .S1(_00450_),
    .X(_04093_));
 sky130_fd_sc_hd__o31a_1 _09704_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[7] ),
    .A2(net3422),
    .A3(_04093_),
    .B1(_00464_),
    .X(_04094_));
 sky130_fd_sc_hd__mux4_1 _09705_ (.A0(_00880_),
    .A1(_03698_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ),
    .X(_04095_));
 sky130_fd_sc_hd__or3_1 _09706_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[7] ),
    .B(_00458_),
    .C(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__mux4_1 _09707_ (.A0(_03484_),
    .A1(_03486_),
    .A2(_03488_),
    .A3(_03490_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ),
    .X(_04097_));
 sky130_fd_sc_hd__mux4_1 _09708_ (.A0(_03806_),
    .A1(_03807_),
    .A2(_03808_),
    .A3(_03809_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ),
    .X(_04098_));
 sky130_fd_sc_hd__mux4_1 _09709_ (.A0(_03493_),
    .A1(_03495_),
    .A2(_03497_),
    .A3(_03499_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ),
    .X(_04099_));
 sky130_fd_sc_hd__and3_1 _09710_ (.A(_00456_),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[8] ),
    .C(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__a31o_1 _09711_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[7] ),
    .A2(_00458_),
    .A3(_04098_),
    .B1(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__a311oi_1 _09712_ (.A1(_00456_),
    .A2(_00458_),
    .A3(_04097_),
    .B1(_04101_),
    .C1(_00464_),
    .Y(_04102_));
 sky130_fd_sc_hd__a31oi_1 _09713_ (.A1(net3423),
    .A2(_04094_),
    .A3(_04096_),
    .B1(_04102_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[1] ));
 sky130_fd_sc_hd__nand3b_2 _09714_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .C(_01415_),
    .Y(_04103_));
 sky130_fd_sc_hd__or3_1 _09715_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_04104_));
 sky130_fd_sc_hd__or2_2 _09716_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__o21a_2 _09717_ (.A1(_04103_),
    .A2(_04105_),
    .B1(_01489_),
    .X(_04106_));
 sky130_fd_sc_hd__mux2_1 _09718_ (.A0(_03865_),
    .A1(net3470),
    .S(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__clkbuf_1 _09719_ (.A(_04107_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _09720_ (.A0(_03872_),
    .A1(net3383),
    .S(_04106_),
    .X(_04108_));
 sky130_fd_sc_hd__clkbuf_1 _09721_ (.A(_04108_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux4_1 _09722_ (.A0(_03478_),
    .A1(_03479_),
    .A2(_03480_),
    .A3(_03481_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[1] ),
    .X(_04109_));
 sky130_fd_sc_hd__inv_2 _09723_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[3] ),
    .Y(_04110_));
 sky130_fd_sc_hd__mux4_1 _09724_ (.A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[1] ),
    .X(_04111_));
 sky130_fd_sc_hd__o21a_1 _09725_ (.A1(_04110_),
    .A2(_04111_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[2] ),
    .X(_04112_));
 sky130_fd_sc_hd__o21ai_1 _09726_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[3] ),
    .A2(_04109_),
    .B1(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__mux4_1 _09727_ (.A0(_03758_),
    .A1(_03759_),
    .A2(_03760_),
    .A3(_03761_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[1] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[0] ),
    .X(_04114_));
 sky130_fd_sc_hd__o31a_1 _09728_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[2] ),
    .A2(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[3] ),
    .A3(_04114_),
    .B1(_00446_),
    .X(_04115_));
 sky130_fd_sc_hd__mux4_1 _09729_ (.A0(_00880_),
    .A1(_03698_),
    .A2(_03473_),
    .A3(_03474_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[1] ),
    .X(_04116_));
 sky130_fd_sc_hd__or3_1 _09730_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[2] ),
    .B(_04110_),
    .C(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__mux4_1 _09731_ (.A0(net21),
    .A1(net22),
    .A2(net23),
    .A3(net24),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[1] ),
    .X(_04118_));
 sky130_fd_sc_hd__inv_2 _09732_ (.A(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__mux4_1 _09733_ (.A0(_03503_),
    .A1(_03504_),
    .A2(_03505_),
    .A3(_03506_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[1] ),
    .X(_04120_));
 sky130_fd_sc_hd__mux4_1 _09734_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[1] ),
    .X(_04121_));
 sky130_fd_sc_hd__and3b_1 _09735_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[2] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[3] ),
    .C(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__a31oi_1 _09736_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[2] ),
    .A2(_04110_),
    .A3(_04120_),
    .B1(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__o311a_1 _09737_ (.A1(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[2] ),
    .A2(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[3] ),
    .A3(_04119_),
    .B1(_04123_),
    .C1(net3743),
    .X(_04124_));
 sky130_fd_sc_hd__a31oi_1 _09738_ (.A1(_04113_),
    .A2(_04115_),
    .A3(_04117_),
    .B1(net3744),
    .Y(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[0] ));
 sky130_fd_sc_hd__mux2_1 _09739_ (.A0(_03874_),
    .A1(net3648),
    .S(_04106_),
    .X(_04125_));
 sky130_fd_sc_hd__clkbuf_1 _09740_ (.A(_04125_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _09741_ (.A0(_03622_),
    .A1(net3509),
    .S(_04106_),
    .X(_04126_));
 sky130_fd_sc_hd__clkbuf_1 _09742_ (.A(_04126_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__clkbuf_2 _09743_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .X(_04127_));
 sky130_fd_sc_hd__inv_2 _09744_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .Y(_04128_));
 sky130_fd_sc_hd__or4_1 _09745_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_04127_),
    .C(_04128_),
    .D(_04103_),
    .X(_04129_));
 sky130_fd_sc_hd__o21a_2 _09746_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .A2(_04129_),
    .B1(_01489_),
    .X(_04130_));
 sky130_fd_sc_hd__mux2_1 _09747_ (.A0(_03865_),
    .A1(net3767),
    .S(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__clkbuf_1 _09748_ (.A(_04131_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _09749_ (.A0(_03872_),
    .A1(net3401),
    .S(_04130_),
    .X(_04132_));
 sky130_fd_sc_hd__clkbuf_1 _09750_ (.A(_04132_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _09751_ (.A0(_03874_),
    .A1(net3399),
    .S(_04130_),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_1 _09752_ (.A(_04133_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _09753_ (.A0(_00192_),
    .A1(net3347),
    .S(_04130_),
    .X(_04134_));
 sky130_fd_sc_hd__clkbuf_1 _09754_ (.A(_04134_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__and3b_2 _09755_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .C(_00311_),
    .X(_04135_));
 sky130_fd_sc_hd__nand2_1 _09756_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_04104_),
    .Y(_04136_));
 sky130_fd_sc_hd__and2_1 _09757_ (.A(_04105_),
    .B(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__inv_2 _09758_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .Y(_04138_));
 sky130_fd_sc_hd__or3_1 _09759_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(_04138_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_04139_));
 sky130_fd_sc_hd__nand2_2 _09760_ (.A(_00170_),
    .B(_04105_),
    .Y(_04140_));
 sky130_fd_sc_hd__nor2_1 _09761_ (.A(_04139_),
    .B(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__inv_2 _09762_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .Y(_04142_));
 sky130_fd_sc_hd__and3b_1 _09763_ (.A_N(_04139_),
    .B(_04142_),
    .C(_04135_),
    .X(_04143_));
 sky130_fd_sc_hd__inv_2 _09764_ (.A(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__a32o_1 _09765_ (.A1(_04135_),
    .A2(_04137_),
    .A3(_04141_),
    .B1(_04144_),
    .B2(net3879),
    .X(_04145_));
 sky130_fd_sc_hd__a21o_1 _09766_ (.A1(_02044_),
    .A2(_04145_),
    .B1(_00210_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__clkinv_2 _09767_ (.A(net3642),
    .Y(_04146_));
 sky130_fd_sc_hd__nand2_1 _09768_ (.A(_01446_),
    .B(_04105_),
    .Y(_04147_));
 sky130_fd_sc_hd__mux2_1 _09769_ (.A0(_04146_),
    .A1(_04147_),
    .S(_04143_),
    .X(_04148_));
 sky130_fd_sc_hd__o21ai_1 _09770_ (.A1(_03914_),
    .A2(_04148_),
    .B1(_03379_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__and2_1 _09771_ (.A(_00187_),
    .B(_04105_),
    .X(_04149_));
 sky130_fd_sc_hd__mux2_1 _09772_ (.A0(net3624),
    .A1(_04149_),
    .S(_04143_),
    .X(_04150_));
 sky130_fd_sc_hd__a21o_1 _09773_ (.A1(_02044_),
    .A2(_04150_),
    .B1(_00262_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__clkinv_2 _09774_ (.A(net3162),
    .Y(_04151_));
 sky130_fd_sc_hd__nand2_2 _09775_ (.A(_01452_),
    .B(_04105_),
    .Y(_04152_));
 sky130_fd_sc_hd__mux2_1 _09776_ (.A0(_04151_),
    .A1(_04152_),
    .S(_04143_),
    .X(_04153_));
 sky130_fd_sc_hd__o21ai_1 _09777_ (.A1(_03914_),
    .A2(_04153_),
    .B1(_03322_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _09778_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(_04103_),
    .Y(_04154_));
 sky130_fd_sc_hd__and3b_2 _09779_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(_04155_));
 sky130_fd_sc_hd__a21oi_4 _09780_ (.A1(_04154_),
    .A2(_04155_),
    .B1(_02686_),
    .Y(_04156_));
 sky130_fd_sc_hd__mux2_1 _09781_ (.A0(_03865_),
    .A1(net3176),
    .S(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__clkbuf_1 _09782_ (.A(_04157_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _09783_ (.A0(_03872_),
    .A1(net3591),
    .S(_04156_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_1 _09784_ (.A(_04158_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _09785_ (.A0(_03874_),
    .A1(net3449),
    .S(_04156_),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_1 _09786_ (.A(_04159_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _09787_ (.A0(_00192_),
    .A1(net3612),
    .S(_04156_),
    .X(_04160_));
 sky130_fd_sc_hd__clkbuf_1 _09788_ (.A(_04160_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4_1 _09789_ (.A(_04127_),
    .B(_04138_),
    .C(_04128_),
    .D(_04154_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_2 _09790_ (.A(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__nand2_1 _09791_ (.A(_04140_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__or2_1 _09792_ (.A(net4182),
    .B(_04162_),
    .X(_04164_));
 sky130_fd_sc_hd__a31o_1 _09793_ (.A1(_03982_),
    .A2(_04163_),
    .A3(_04164_),
    .B1(_03316_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _09794_ (.A(_04147_),
    .B(_04162_),
    .Y(_04165_));
 sky130_fd_sc_hd__or2_1 _09795_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ),
    .B(_04162_),
    .X(_04166_));
 sky130_fd_sc_hd__a31o_1 _09796_ (.A1(_03982_),
    .A2(_04165_),
    .A3(_04166_),
    .B1(_01772_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__or2b_1 _09797_ (.A(_04149_),
    .B_N(_04162_),
    .X(_04167_));
 sky130_fd_sc_hd__or2_1 _09798_ (.A(net4111),
    .B(_04162_),
    .X(_04168_));
 sky130_fd_sc_hd__a31o_1 _09799_ (.A1(_03982_),
    .A2(_04167_),
    .A3(_04168_),
    .B1(_01851_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _09800_ (.A(net3930),
    .B(_04162_),
    .Y(_04169_));
 sky130_fd_sc_hd__a211o_1 _09801_ (.A1(_04152_),
    .A2(_04162_),
    .B1(_04169_),
    .C1(_00228_),
    .X(_04170_));
 sky130_fd_sc_hd__nand2_1 _09802_ (.A(_03166_),
    .B(_04170_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _09803_ (.A1(_04127_),
    .A2(_04138_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .A4(_04154_),
    .B1(_00249_),
    .X(_04171_));
 sky130_fd_sc_hd__mux2_1 _09804_ (.A0(net4100),
    .A1(_00235_),
    .S(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _09805_ (.A(_04172_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _09806_ (.A0(net3894),
    .A1(_00292_),
    .S(_04171_),
    .X(_04173_));
 sky130_fd_sc_hd__clkbuf_1 _09807_ (.A(_04173_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _09808_ (.A0(net3779),
    .A1(_00188_),
    .S(_04171_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _09809_ (.A(_04174_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _09810_ (.A0(net3825),
    .A1(_00527_),
    .S(_04171_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _09811_ (.A(_04175_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4_2 _09812_ (.A(_04127_),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .C(_04128_),
    .D(_04154_),
    .X(_04176_));
 sky130_fd_sc_hd__or2_1 _09813_ (.A(net4167),
    .B(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__nand2_1 _09814_ (.A(_04140_),
    .B(_04176_),
    .Y(_04178_));
 sky130_fd_sc_hd__a31o_1 _09815_ (.A1(_03982_),
    .A2(_04177_),
    .A3(_04178_),
    .B1(_01766_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _09816_ (.A0(_00984_),
    .A1(_04147_),
    .S(_04176_),
    .X(_04179_));
 sky130_fd_sc_hd__o21ai_1 _09817_ (.A1(_03914_),
    .A2(_04179_),
    .B1(_03379_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _09818_ (.A0(net4190),
    .A1(_04149_),
    .S(_04176_),
    .X(_04180_));
 sky130_fd_sc_hd__a21o_1 _09819_ (.A1(_00223_),
    .A2(_04180_),
    .B1(_00262_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__clkbuf_4 _09820_ (.A(_01764_),
    .X(_04181_));
 sky130_fd_sc_hd__mux2_1 _09821_ (.A0(_00994_),
    .A1(_04152_),
    .S(_04176_),
    .X(_04182_));
 sky130_fd_sc_hd__o21ai_1 _09822_ (.A1(_04181_),
    .A2(_04182_),
    .B1(_03322_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _09823_ (.A1(_04127_),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .A4(_04154_),
    .B1(_00249_),
    .X(_04183_));
 sky130_fd_sc_hd__mux2_1 _09824_ (.A0(net4055),
    .A1(_00235_),
    .S(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_1 _09825_ (.A(_04184_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _09826_ (.A0(net4194),
    .A1(_00292_),
    .S(_04183_),
    .X(_04185_));
 sky130_fd_sc_hd__clkbuf_1 _09827_ (.A(_04185_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _09828_ (.A0(net3674),
    .A1(_00188_),
    .S(_04183_),
    .X(_04186_));
 sky130_fd_sc_hd__clkbuf_1 _09829_ (.A(_04186_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _09830_ (.A0(net3971),
    .A1(_00527_),
    .S(_04183_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _09831_ (.A(_04187_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__o31a_2 _09832_ (.A1(_04142_),
    .A2(_04103_),
    .A3(_04104_),
    .B1(_02847_),
    .X(_04188_));
 sky130_fd_sc_hd__mux2_1 _09833_ (.A0(_03865_),
    .A1(net3974),
    .S(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _09834_ (.A(_04189_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _09835_ (.A0(_03872_),
    .A1(net3630),
    .S(_04188_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _09836_ (.A(_04190_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _09837_ (.A0(_03874_),
    .A1(net3647),
    .S(_04188_),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _09838_ (.A(_04191_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _09839_ (.A0(_00192_),
    .A1(net3904),
    .S(_04188_),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _09840_ (.A(_04192_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _09841_ (.A(_04103_),
    .B(_04137_),
    .X(_04193_));
 sky130_fd_sc_hd__o41a_2 _09842_ (.A1(_04127_),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .A3(_04128_),
    .A4(_04193_),
    .B1(_00407_),
    .X(_04194_));
 sky130_fd_sc_hd__mux2_1 _09843_ (.A0(_03865_),
    .A1(net3626),
    .S(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _09844_ (.A(_04195_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _09845_ (.A0(_03872_),
    .A1(net3468),
    .S(_04194_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _09846_ (.A(_04196_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _09847_ (.A0(_03874_),
    .A1(net3241),
    .S(_04194_),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_1 _09848_ (.A(_04197_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _09849_ (.A0(_00192_),
    .A1(net3477),
    .S(_04194_),
    .X(_04198_));
 sky130_fd_sc_hd__clkbuf_1 _09850_ (.A(_04198_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _09851_ (.A(_04139_),
    .B(_04193_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand2_1 _09852_ (.A(_04140_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__or2_1 _09853_ (.A(net4075),
    .B(_04199_),
    .X(_04201_));
 sky130_fd_sc_hd__a31o_1 _09854_ (.A1(_03982_),
    .A2(_04200_),
    .A3(_04201_),
    .B1(_01766_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__or2_1 _09855_ (.A(net3928),
    .B(_04199_),
    .X(_04202_));
 sky130_fd_sc_hd__nand2_1 _09856_ (.A(_04147_),
    .B(_04199_),
    .Y(_04203_));
 sky130_fd_sc_hd__a31o_1 _09857_ (.A1(_03982_),
    .A2(_04202_),
    .A3(_04203_),
    .B1(_01772_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__mux2_1 _09858_ (.A0(net3337),
    .A1(_04149_),
    .S(_04199_),
    .X(_04204_));
 sky130_fd_sc_hd__a21o_1 _09859_ (.A1(_00223_),
    .A2(_04204_),
    .B1(_00262_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__nor2_1 _09860_ (.A(net3983),
    .B(_04199_),
    .Y(_04205_));
 sky130_fd_sc_hd__a211o_1 _09861_ (.A1(_04152_),
    .A2(_04199_),
    .B1(_04205_),
    .C1(_00228_),
    .X(_04206_));
 sky130_fd_sc_hd__nand2_1 _09862_ (.A(_00276_),
    .B(_04206_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3b_1 _09863_ (.A_N(_04137_),
    .B(_04155_),
    .C(_04135_),
    .X(_04207_));
 sky130_fd_sc_hd__a31oi_4 _09864_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .A2(_04135_),
    .A3(_04155_),
    .B1(_02637_),
    .Y(_04208_));
 sky130_fd_sc_hd__a221o_1 _09865_ (.A1(_00288_),
    .A2(_04207_),
    .B1(_04208_),
    .B2(net3166),
    .C1(_00209_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _09866_ (.A1(_00293_),
    .A2(_04207_),
    .B1(_04208_),
    .B2(net3218),
    .C1(_02872_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _09867_ (.A1(_00295_),
    .A2(_04207_),
    .B1(_04208_),
    .B2(net3203),
    .C1(_00221_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__nor2_1 _09868_ (.A(_02759_),
    .B(_01054_),
    .Y(_04209_));
 sky130_fd_sc_hd__mux2_1 _09869_ (.A0(_03992_),
    .A1(_04209_),
    .S(_03993_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _09870_ (.A(_04210_),
    .X(_00002_));
 sky130_fd_sc_hd__mux4_1 _09871_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ),
    .X(_04211_));
 sky130_fd_sc_hd__mux4_1 _09872_ (.A0(_03816_),
    .A1(_03817_),
    .A2(_03818_),
    .A3(_03819_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ),
    .X(_04212_));
 sky130_fd_sc_hd__or2_1 _09873_ (.A(_00653_),
    .B(_04212_),
    .X(_04213_));
 sky130_fd_sc_hd__o211a_1 _09874_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[38] ),
    .A2(_04211_),
    .B1(_04213_),
    .C1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[37] ),
    .X(_04214_));
 sky130_fd_sc_hd__buf_2 _09875_ (.A(_01580_),
    .X(_04215_));
 sky130_fd_sc_hd__buf_2 _09876_ (.A(_01673_),
    .X(_04216_));
 sky130_fd_sc_hd__buf_2 _09877_ (.A(_01759_),
    .X(_04217_));
 sky130_fd_sc_hd__buf_2 _09878_ (.A(_01849_),
    .X(_04218_));
 sky130_fd_sc_hd__mux4_1 _09879_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04217_),
    .A3(_04218_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ),
    .X(_04219_));
 sky130_fd_sc_hd__nor3_1 _09880_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[37] ),
    .B(_00653_),
    .C(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__nor2_1 _09881_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[37] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[38] ),
    .Y(_04221_));
 sky130_fd_sc_hd__mux4_1 _09882_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .S0(_00649_),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ),
    .X(_04222_));
 sky130_fd_sc_hd__a21o_1 _09883_ (.A1(_04221_),
    .A2(_04222_),
    .B1(net3307),
    .X(_04223_));
 sky130_fd_sc_hd__mux4_1 _09884_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ),
    .X(_04224_));
 sky130_fd_sc_hd__mux4_1 _09885_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ),
    .X(_04225_));
 sky130_fd_sc_hd__mux4_1 _09886_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ),
    .X(_04226_));
 sky130_fd_sc_hd__and3_1 _09887_ (.A(_00651_),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[38] ),
    .C(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__a31o_1 _09888_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[37] ),
    .A2(_00653_),
    .A3(_04225_),
    .B1(_04227_),
    .X(_04228_));
 sky130_fd_sc_hd__a211o_1 _09889_ (.A1(_04221_),
    .A2(_04224_),
    .B1(_04228_),
    .C1(_00655_),
    .X(_04229_));
 sky130_fd_sc_hd__o31a_1 _09890_ (.A1(_04214_),
    .A2(_04220_),
    .A3(_04223_),
    .B1(_04229_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[7] ));
 sky130_fd_sc_hd__mux4_1 _09891_ (.A0(_03478_),
    .A1(_03479_),
    .A2(_03480_),
    .A3(_03481_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ),
    .X(_04230_));
 sky130_fd_sc_hd__inv_2 _09892_ (.A(net3826),
    .Y(_04231_));
 sky130_fd_sc_hd__mux4_1 _09893_ (.A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ),
    .X(_04232_));
 sky130_fd_sc_hd__o21a_1 _09894_ (.A1(_04231_),
    .A2(_04232_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ),
    .X(_04233_));
 sky130_fd_sc_hd__o21ai_1 _09895_ (.A1(net3826),
    .A2(_04230_),
    .B1(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__mux4_1 _09896_ (.A0(_03760_),
    .A1(_03761_),
    .A2(_03758_),
    .A3(_03759_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ),
    .S1(_00636_),
    .X(_04235_));
 sky130_fd_sc_hd__inv_2 _09897_ (.A(net3724),
    .Y(_04236_));
 sky130_fd_sc_hd__o31a_1 _09898_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ),
    .A2(net3826),
    .A3(_04235_),
    .B1(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__mux4_1 _09899_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ),
    .X(_04238_));
 sky130_fd_sc_hd__or3_1 _09900_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ),
    .B(_04231_),
    .C(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__mux4_1 _09901_ (.A0(net25),
    .A1(net26),
    .A2(net12),
    .A3(net13),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ),
    .X(_04240_));
 sky130_fd_sc_hd__a31o_1 _09902_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ),
    .A2(_04231_),
    .A3(_04240_),
    .B1(_04236_),
    .X(_04241_));
 sky130_fd_sc_hd__mux4_1 _09903_ (.A0(_03546_),
    .A1(_03547_),
    .A2(_03548_),
    .A3(_03549_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ),
    .X(_04242_));
 sky130_fd_sc_hd__or3b_1 _09904_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ),
    .B(_04231_),
    .C_N(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__mux4_1 _09905_ (.A0(net21),
    .A1(net22),
    .A2(net23),
    .A3(net24),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ),
    .X(_04244_));
 sky130_fd_sc_hd__or3b_1 _09906_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[33] ),
    .C_N(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__and3b_1 _09907_ (.A_N(_04241_),
    .B(_04243_),
    .C(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__a31oi_1 _09908_ (.A1(net3827),
    .A2(_04237_),
    .A3(_04239_),
    .B1(_04246_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[6] ));
 sky130_fd_sc_hd__mux4_1 _09909_ (.A0(_03478_),
    .A1(_03479_),
    .A2(_03480_),
    .A3(_03481_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ),
    .X(_04247_));
 sky130_fd_sc_hd__mux4_1 _09910_ (.A0(_03516_),
    .A1(_03517_),
    .A2(_03518_),
    .A3(_03519_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ),
    .X(_04248_));
 sky130_fd_sc_hd__o21a_1 _09911_ (.A1(_00631_),
    .A2(_04248_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[27] ),
    .X(_04249_));
 sky130_fd_sc_hd__o21ai_1 _09912_ (.A1(net3738),
    .A2(_04247_),
    .B1(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__mux4_1 _09913_ (.A0(_03760_),
    .A1(_03761_),
    .A2(_03758_),
    .A3(_03759_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ),
    .S1(_00625_),
    .X(_04251_));
 sky130_fd_sc_hd__o31a_1 _09914_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[27] ),
    .A2(net3738),
    .A3(_04251_),
    .B1(_00634_),
    .X(_04252_));
 sky130_fd_sc_hd__mux4_1 _09915_ (.A0(_01580_),
    .A1(_01673_),
    .A2(_01759_),
    .A3(_01849_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ),
    .X(_04253_));
 sky130_fd_sc_hd__or3_1 _09916_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[27] ),
    .B(_00631_),
    .C(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__mux4_1 _09917_ (.A0(_03484_),
    .A1(_03486_),
    .A2(_03488_),
    .A3(_03490_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ),
    .X(_04255_));
 sky130_fd_sc_hd__mux4_1 _09918_ (.A0(_03806_),
    .A1(_03807_),
    .A2(_03808_),
    .A3(_03809_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ),
    .X(_04256_));
 sky130_fd_sc_hd__mux4_1 _09919_ (.A0(_03493_),
    .A1(_03495_),
    .A2(_03497_),
    .A3(_03499_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[25] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ),
    .X(_04257_));
 sky130_fd_sc_hd__and3_1 _09920_ (.A(_00629_),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[28] ),
    .C(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__a31o_1 _09921_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[27] ),
    .A2(_00631_),
    .A3(_04256_),
    .B1(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__a311oi_1 _09922_ (.A1(_00629_),
    .A2(_00631_),
    .A3(_04255_),
    .B1(_04259_),
    .C1(_00634_),
    .Y(_04260_));
 sky130_fd_sc_hd__a31oi_1 _09923_ (.A1(net3739),
    .A2(_04252_),
    .A3(_04254_),
    .B1(_04260_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[5] ));
 sky130_fd_sc_hd__mux4_1 _09924_ (.A0(_02226_),
    .A1(_02320_),
    .A2(_02408_),
    .A3(_02491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ),
    .X(_04261_));
 sky130_fd_sc_hd__mux4_1 _09925_ (.A0(net11),
    .A1(net18),
    .A2(net19),
    .A3(net20),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ),
    .X(_04262_));
 sky130_fd_sc_hd__or2_1 _09926_ (.A(_00619_),
    .B(_04262_),
    .X(_04263_));
 sky130_fd_sc_hd__o211a_1 _09927_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[23] ),
    .A2(_04261_),
    .B1(_04263_),
    .C1(net3282),
    .X(_04264_));
 sky130_fd_sc_hd__mux4_1 _09928_ (.A0(_03780_),
    .A1(_03781_),
    .A2(_03782_),
    .A3(_03783_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ),
    .S1(_00610_),
    .X(_04265_));
 sky130_fd_sc_hd__and3_1 _09929_ (.A(_00617_),
    .B(_00619_),
    .C(_04265_),
    .X(_04266_));
 sky130_fd_sc_hd__mux4_1 _09930_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04217_),
    .A3(_04218_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ),
    .X(_04267_));
 sky130_fd_sc_hd__nor3_1 _09931_ (.A(net3282),
    .B(_00619_),
    .C(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__mux4_1 _09932_ (.A0(_03484_),
    .A1(_03486_),
    .A2(_03488_),
    .A3(_03490_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ),
    .X(_04269_));
 sky130_fd_sc_hd__mux4_1 _09933_ (.A0(_03806_),
    .A1(_03807_),
    .A2(_03808_),
    .A3(_03809_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ),
    .X(_04270_));
 sky130_fd_sc_hd__mux4_1 _09934_ (.A0(net14),
    .A1(net15),
    .A2(net16),
    .A3(net17),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ),
    .X(_04271_));
 sky130_fd_sc_hd__and3_1 _09935_ (.A(_00617_),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[23] ),
    .C(_04271_),
    .X(_04272_));
 sky130_fd_sc_hd__a31o_1 _09936_ (.A1(net3282),
    .A2(_00619_),
    .A3(_04270_),
    .B1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__a311o_1 _09937_ (.A1(_00617_),
    .A2(_00619_),
    .A3(_04269_),
    .B1(_04273_),
    .C1(_00622_),
    .X(_04274_));
 sky130_fd_sc_hd__o41a_1 _09938_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[24] ),
    .A2(net3283),
    .A3(_04266_),
    .A4(_04268_),
    .B1(_04274_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[4] ));
 sky130_fd_sc_hd__mux4_1 _09939_ (.A0(_02226_),
    .A1(_02320_),
    .A2(_02408_),
    .A3(_02491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ),
    .X(_04275_));
 sky130_fd_sc_hd__inv_2 _09940_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ),
    .Y(_04276_));
 sky130_fd_sc_hd__mux4_1 _09941_ (.A0(_03816_),
    .A1(_03817_),
    .A2(_03818_),
    .A3(_03819_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ),
    .X(_04277_));
 sky130_fd_sc_hd__or2_1 _09942_ (.A(_04276_),
    .B(_04277_),
    .X(_04278_));
 sky130_fd_sc_hd__o211a_1 _09943_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ),
    .A2(_04275_),
    .B1(_04278_),
    .C1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ),
    .X(_04279_));
 sky130_fd_sc_hd__mux4_1 _09944_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04217_),
    .A3(_04218_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ),
    .X(_04280_));
 sky130_fd_sc_hd__nor3_1 _09945_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ),
    .B(_04276_),
    .C(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__nor2_1 _09946_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ),
    .Y(_04282_));
 sky130_fd_sc_hd__mux4_1 _09947_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ),
    .S1(_00597_),
    .X(_04283_));
 sky130_fd_sc_hd__a21o_1 _09948_ (.A1(_04282_),
    .A2(_04283_),
    .B1(net3890),
    .X(_04284_));
 sky130_fd_sc_hd__mux4_1 _09949_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ),
    .X(_04285_));
 sky130_fd_sc_hd__mux4_1 _09950_ (.A0(_03541_),
    .A1(_03542_),
    .A2(_03543_),
    .A3(_03544_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ),
    .X(_04286_));
 sky130_fd_sc_hd__mux4_1 _09951_ (.A0(_03493_),
    .A1(_03495_),
    .A2(_03497_),
    .A3(_03499_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[15] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ),
    .X(_04287_));
 sky130_fd_sc_hd__and3b_1 _09952_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ),
    .C(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__a31o_1 _09953_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ),
    .A2(_04276_),
    .A3(_04286_),
    .B1(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__inv_2 _09954_ (.A(net3890),
    .Y(_04290_));
 sky130_fd_sc_hd__a211o_1 _09955_ (.A1(_04282_),
    .A2(_04285_),
    .B1(_04289_),
    .C1(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__o31a_1 _09956_ (.A1(_04279_),
    .A2(_04281_),
    .A3(_04284_),
    .B1(_04291_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[3] ));
 sky130_fd_sc_hd__mux4_1 _09957_ (.A0(_03478_),
    .A1(_03479_),
    .A2(_03480_),
    .A3(_03481_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[11] ),
    .X(_04292_));
 sky130_fd_sc_hd__mux4_1 _09958_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[11] ),
    .X(_04293_));
 sky130_fd_sc_hd__o21a_1 _09959_ (.A1(_00592_),
    .A2(_04293_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[12] ),
    .X(_04294_));
 sky130_fd_sc_hd__o21ai_1 _09960_ (.A1(net3946),
    .A2(_04292_),
    .B1(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__mux4_1 _09961_ (.A0(_03760_),
    .A1(_03761_),
    .A2(_03758_),
    .A3(_03759_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[11] ),
    .S1(_00584_),
    .X(_04296_));
 sky130_fd_sc_hd__o31a_1 _09962_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[12] ),
    .A2(net3946),
    .A3(_04296_),
    .B1(_00594_),
    .X(_04297_));
 sky130_fd_sc_hd__mux4_1 _09963_ (.A0(_01580_),
    .A1(_01673_),
    .A2(_01759_),
    .A3(_01849_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[11] ),
    .X(_04298_));
 sky130_fd_sc_hd__or3_1 _09964_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[12] ),
    .B(_00592_),
    .C(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__mux4_1 _09965_ (.A0(_03484_),
    .A1(_03486_),
    .A2(_03488_),
    .A3(_03490_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[11] ),
    .X(_04300_));
 sky130_fd_sc_hd__mux4_1 _09966_ (.A0(_03806_),
    .A1(_03807_),
    .A2(_03808_),
    .A3(_03809_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[11] ),
    .X(_04301_));
 sky130_fd_sc_hd__mux4_1 _09967_ (.A0(net14),
    .A1(net15),
    .A2(net16),
    .A3(net17),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[10] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[11] ),
    .X(_04302_));
 sky130_fd_sc_hd__and3_1 _09968_ (.A(_00588_),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[13] ),
    .C(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__a31o_1 _09969_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[12] ),
    .A2(_00592_),
    .A3(_04301_),
    .B1(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__a311oi_1 _09970_ (.A1(_00588_),
    .A2(_00592_),
    .A3(_04300_),
    .B1(_04304_),
    .C1(_00594_),
    .Y(_04305_));
 sky130_fd_sc_hd__a31oi_1 _09971_ (.A1(net3947),
    .A2(_04297_),
    .A3(_04299_),
    .B1(_04305_),
    .Y(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[2] ));
 sky130_fd_sc_hd__mux4_1 _09972_ (.A0(_02226_),
    .A1(_02320_),
    .A2(_02408_),
    .A3(_02491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ),
    .X(_04306_));
 sky130_fd_sc_hd__mux4_1 _09973_ (.A0(net11),
    .A1(net18),
    .A2(net19),
    .A3(net20),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ),
    .X(_04307_));
 sky130_fd_sc_hd__or2_1 _09974_ (.A(_00577_),
    .B(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__o211a_1 _09975_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[8] ),
    .A2(_04306_),
    .B1(_04308_),
    .C1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[7] ),
    .X(_04309_));
 sky130_fd_sc_hd__mux4_1 _09976_ (.A0(_00785_),
    .A1(_01144_),
    .A2(_01228_),
    .A3(_01057_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ),
    .S1(_00569_),
    .X(_04310_));
 sky130_fd_sc_hd__and3_1 _09977_ (.A(_00575_),
    .B(_00577_),
    .C(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__mux4_1 _09978_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04217_),
    .A3(_04218_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ),
    .X(_04312_));
 sky130_fd_sc_hd__nor3_1 _09979_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[7] ),
    .B(_00577_),
    .C(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__mux4_1 _09980_ (.A0(_03484_),
    .A1(_03486_),
    .A2(_03488_),
    .A3(_03490_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ),
    .X(_04314_));
 sky130_fd_sc_hd__mux4_1 _09981_ (.A0(_03806_),
    .A1(_03807_),
    .A2(_03808_),
    .A3(_03809_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ),
    .X(_04315_));
 sky130_fd_sc_hd__mux4_1 _09982_ (.A0(net14),
    .A1(net15),
    .A2(net16),
    .A3(net17),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ),
    .X(_04316_));
 sky130_fd_sc_hd__and3_1 _09983_ (.A(_00575_),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[8] ),
    .C(_04316_),
    .X(_04317_));
 sky130_fd_sc_hd__a31o_1 _09984_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[7] ),
    .A2(_00577_),
    .A3(_04315_),
    .B1(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__a311o_1 _09985_ (.A1(_00575_),
    .A2(_00577_),
    .A3(_04314_),
    .B1(_04318_),
    .C1(_00582_),
    .X(_04319_));
 sky130_fd_sc_hd__o41a_1 _09986_ (.A1(net3287),
    .A2(_04309_),
    .A3(_04311_),
    .A4(_04313_),
    .B1(_04319_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[1] ));
 sky130_fd_sc_hd__mux4_1 _09987_ (.A0(_02226_),
    .A1(_02320_),
    .A2(_02408_),
    .A3(_02491_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ),
    .X(_04320_));
 sky130_fd_sc_hd__inv_2 _09988_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ),
    .Y(_04321_));
 sky130_fd_sc_hd__mux4_1 _09989_ (.A0(_03816_),
    .A1(_03817_),
    .A2(_03818_),
    .A3(_03819_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ),
    .X(_04322_));
 sky130_fd_sc_hd__or2_1 _09990_ (.A(_04321_),
    .B(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__o211a_1 _09991_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ),
    .A2(_04320_),
    .B1(_04323_),
    .C1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ),
    .X(_04324_));
 sky130_fd_sc_hd__mux4_1 _09992_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04217_),
    .A3(_04218_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ),
    .X(_04325_));
 sky130_fd_sc_hd__nor3_1 _09993_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ),
    .B(_04321_),
    .C(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__nor2_1 _09994_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ),
    .Y(_04327_));
 sky130_fd_sc_hd__mux4_1 _09995_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ),
    .X(_04328_));
 sky130_fd_sc_hd__a21o_1 _09996_ (.A1(_04327_),
    .A2(_04328_),
    .B1(net3688),
    .X(_04329_));
 sky130_fd_sc_hd__mux4_1 _09997_ (.A0(_03536_),
    .A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ),
    .X(_04330_));
 sky130_fd_sc_hd__mux4_1 _09998_ (.A0(_03806_),
    .A1(_03807_),
    .A2(_03808_),
    .A3(_03809_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ),
    .X(_04331_));
 sky130_fd_sc_hd__mux4_1 _09999_ (.A0(_03493_),
    .A1(_03495_),
    .A2(_03497_),
    .A3(_03499_),
    .S0(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ),
    .X(_04332_));
 sky130_fd_sc_hd__and3b_1 _10000_ (.A_N(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ),
    .C(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__a31o_1 _10001_ (.A1(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ),
    .A2(_04321_),
    .A3(_04331_),
    .B1(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__a211o_1 _10002_ (.A1(_04327_),
    .A2(_04330_),
    .B1(_04334_),
    .C1(_00565_),
    .X(_04335_));
 sky130_fd_sc_hd__o31a_1 _10003_ (.A1(_04324_),
    .A2(_04326_),
    .A3(_04329_),
    .B1(_04335_),
    .X(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[0] ));
 sky130_fd_sc_hd__nand3b_2 _10004_ (.A_N(\c.genblk1.genblk1.subs.c0.cfgd ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .C(_01878_),
    .Y(_04336_));
 sky130_fd_sc_hd__or3_1 _10005_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_04337_));
 sky130_fd_sc_hd__or2_1 _10006_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10007_ (.A(_04338_),
    .X(_04339_));
 sky130_fd_sc_hd__o21a_2 _10008_ (.A1(_04336_),
    .A2(_04339_),
    .B1(_01489_),
    .X(_04340_));
 sky130_fd_sc_hd__mux2_1 _10009_ (.A0(_00172_),
    .A1(net3300),
    .S(_04340_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_1 _10010_ (.A(_04341_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ));
 sky130_fd_sc_hd__mux2_1 _10011_ (.A0(_00185_),
    .A1(net3606),
    .S(_04340_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _10012_ (.A(_04342_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ));
 sky130_fd_sc_hd__mux2_1 _10013_ (.A0(_00189_),
    .A1(net3329),
    .S(_04340_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _10014_ (.A(_04343_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ));
 sky130_fd_sc_hd__mux2_1 _10015_ (.A0(_00192_),
    .A1(net3651),
    .S(_04340_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _10016_ (.A(_04344_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ));
 sky130_fd_sc_hd__clkbuf_2 _10017_ (.A(net4001),
    .X(_04345_));
 sky130_fd_sc_hd__or3b_1 _10018_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .B(_04345_),
    .C_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_04346_));
 sky130_fd_sc_hd__o31a_2 _10019_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .A2(_04336_),
    .A3(_04346_),
    .B1(_02847_),
    .X(_04347_));
 sky130_fd_sc_hd__mux2_1 _10020_ (.A0(_00172_),
    .A1(net3410),
    .S(_04347_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _10021_ (.A(_04348_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ));
 sky130_fd_sc_hd__mux2_1 _10022_ (.A0(_00185_),
    .A1(net3302),
    .S(_04347_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _10023_ (.A(_04349_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ));
 sky130_fd_sc_hd__mux2_1 _10024_ (.A0(_00189_),
    .A1(net3364),
    .S(_04347_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_1 _10025_ (.A(_04350_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ));
 sky130_fd_sc_hd__mux2_1 _10026_ (.A0(_00192_),
    .A1(net3421),
    .S(_04347_),
    .X(_04351_));
 sky130_fd_sc_hd__clkbuf_1 _10027_ (.A(_04351_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ));
 sky130_fd_sc_hd__inv_2 _10028_ (.A(_04345_),
    .Y(_04352_));
 sky130_fd_sc_hd__or3_2 _10029_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .B(_04352_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_04353_));
 sky130_fd_sc_hd__and3b_1 _10030_ (.A_N(\c.genblk1.genblk1.subs.c0.cfgd ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .C(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ),
    .X(_04354_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10031_ (.A(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__nand2_1 _10032_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_04337_),
    .Y(_04356_));
 sky130_fd_sc_hd__and2_1 _10033_ (.A(_04339_),
    .B(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__nand2_1 _10034_ (.A(_04355_),
    .B(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__nand2_1 _10035_ (.A(_02003_),
    .B(_04339_),
    .Y(_04359_));
 sky130_fd_sc_hd__or3_1 _10036_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_04336_),
    .C(_04353_),
    .X(_04360_));
 sky130_fd_sc_hd__nand2_1 _10037_ (.A(net3835),
    .B(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__o31a_1 _10038_ (.A1(_04353_),
    .A2(_04358_),
    .A3(_04359_),
    .B1(_04361_),
    .X(_04362_));
 sky130_fd_sc_hd__o21ai_1 _10039_ (.A1(_04181_),
    .A2(_04362_),
    .B1(_00237_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ));
 sky130_fd_sc_hd__nand2_1 _10040_ (.A(_01446_),
    .B(_04339_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand2_1 _10041_ (.A(net3789),
    .B(_04360_),
    .Y(_04364_));
 sky130_fd_sc_hd__o31a_1 _10042_ (.A1(_04353_),
    .A2(_04358_),
    .A3(_04363_),
    .B1(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__o21ai_1 _10043_ (.A1(_04181_),
    .A2(_04365_),
    .B1(_03379_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ));
 sky130_fd_sc_hd__nand2_1 _10044_ (.A(_02573_),
    .B(_04339_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand2_1 _10045_ (.A(net3229),
    .B(_04360_),
    .Y(_04367_));
 sky130_fd_sc_hd__o31a_1 _10046_ (.A1(_04353_),
    .A2(_04358_),
    .A3(_04366_),
    .B1(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__o21ai_1 _10047_ (.A1(_04181_),
    .A2(_04368_),
    .B1(_00251_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ));
 sky130_fd_sc_hd__nand2_1 _10048_ (.A(_00264_),
    .B(_04339_),
    .Y(_04369_));
 sky130_fd_sc_hd__nand2_1 _10049_ (.A(net3221),
    .B(_04360_),
    .Y(_04370_));
 sky130_fd_sc_hd__o31a_1 _10050_ (.A1(_04353_),
    .A2(_04358_),
    .A3(_04369_),
    .B1(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__o21ai_1 _10051_ (.A1(_04181_),
    .A2(_04371_),
    .B1(_03322_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ));
 sky130_fd_sc_hd__nor2_2 _10052_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_04336_),
    .Y(_04372_));
 sky130_fd_sc_hd__and3b_1 _10053_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .B(_04345_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(_04373_));
 sky130_fd_sc_hd__a21oi_4 _10054_ (.A1(_04372_),
    .A2(_04373_),
    .B1(_00181_),
    .Y(_04374_));
 sky130_fd_sc_hd__mux2_1 _10055_ (.A0(_00172_),
    .A1(net3385),
    .S(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_1 _10056_ (.A(_04375_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ));
 sky130_fd_sc_hd__mux2_1 _10057_ (.A0(_00185_),
    .A1(net3559),
    .S(_04374_),
    .X(_04376_));
 sky130_fd_sc_hd__clkbuf_1 _10058_ (.A(_04376_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ));
 sky130_fd_sc_hd__mux2_1 _10059_ (.A0(_00189_),
    .A1(net3594),
    .S(_04374_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_1 _10060_ (.A(_04377_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ));
 sky130_fd_sc_hd__mux2_1 _10061_ (.A0(_00192_),
    .A1(net3370),
    .S(_04374_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_1 _10062_ (.A(_04378_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ));
 sky130_fd_sc_hd__and4bb_2 _10063_ (.A_N(_04345_),
    .B_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .C(_04372_),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .X(_04379_));
 sky130_fd_sc_hd__nand2_1 _10064_ (.A(_04359_),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__or2_1 _10065_ (.A(net4155),
    .B(_04379_),
    .X(_04381_));
 sky130_fd_sc_hd__a31o_1 _10066_ (.A1(_03982_),
    .A2(_04380_),
    .A3(_04381_),
    .B1(_01766_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ));
 sky130_fd_sc_hd__nand2_1 _10067_ (.A(_04363_),
    .B(_04379_),
    .Y(_04382_));
 sky130_fd_sc_hd__or2_1 _10068_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .B(_04379_),
    .X(_04383_));
 sky130_fd_sc_hd__a31o_1 _10069_ (.A1(_03982_),
    .A2(_04382_),
    .A3(_04383_),
    .B1(_01772_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ));
 sky130_fd_sc_hd__nand2_1 _10070_ (.A(_04366_),
    .B(_04379_),
    .Y(_04384_));
 sky130_fd_sc_hd__or2_1 _10071_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .B(_04379_),
    .X(_04385_));
 sky130_fd_sc_hd__a31o_1 _10072_ (.A1(_03982_),
    .A2(_04384_),
    .A3(_04385_),
    .B1(_01851_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ));
 sky130_fd_sc_hd__nor2_1 _10073_ (.A(net4029),
    .B(_04379_),
    .Y(_04386_));
 sky130_fd_sc_hd__a211o_1 _10074_ (.A1(_04369_),
    .A2(_04379_),
    .B1(_04386_),
    .C1(_00228_),
    .X(_04387_));
 sky130_fd_sc_hd__nand2_1 _10075_ (.A(_00276_),
    .B(_04387_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ));
 sky130_fd_sc_hd__a41o_2 _10076_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .A2(_04352_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .A4(_04372_),
    .B1(_00249_),
    .X(_04388_));
 sky130_fd_sc_hd__mux2_1 _10077_ (.A0(net4002),
    .A1(_00235_),
    .S(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__clkbuf_1 _10078_ (.A(_04389_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ));
 sky130_fd_sc_hd__mux2_1 _10079_ (.A0(net4152),
    .A1(_00292_),
    .S(_04388_),
    .X(_04390_));
 sky130_fd_sc_hd__clkbuf_1 _10080_ (.A(_04390_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ));
 sky130_fd_sc_hd__mux2_1 _10081_ (.A0(net4026),
    .A1(_00188_),
    .S(_04388_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _10082_ (.A(_04391_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ));
 sky130_fd_sc_hd__mux2_1 _10083_ (.A0(net3669),
    .A1(_00527_),
    .S(_04388_),
    .X(_04392_));
 sky130_fd_sc_hd__clkbuf_1 _10084_ (.A(_04392_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ));
 sky130_fd_sc_hd__and4b_2 _10085_ (.A_N(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .B(_04372_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .D(_04345_),
    .X(_04393_));
 sky130_fd_sc_hd__mux2_1 _10086_ (.A0(_01075_),
    .A1(_04359_),
    .S(_04393_),
    .X(_04394_));
 sky130_fd_sc_hd__o21ai_1 _10087_ (.A1(_04181_),
    .A2(_04394_),
    .B1(_00237_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ));
 sky130_fd_sc_hd__mux2_1 _10088_ (.A0(_01078_),
    .A1(_04363_),
    .S(_04393_),
    .X(_04395_));
 sky130_fd_sc_hd__o21ai_1 _10089_ (.A1(_04181_),
    .A2(_04395_),
    .B1(_00305_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ));
 sky130_fd_sc_hd__mux2_1 _10090_ (.A0(_01080_),
    .A1(_04366_),
    .S(_04393_),
    .X(_04396_));
 sky130_fd_sc_hd__o21ai_1 _10091_ (.A1(_04181_),
    .A2(_04396_),
    .B1(_00251_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ));
 sky130_fd_sc_hd__mux2_1 _10092_ (.A0(_01070_),
    .A1(_04369_),
    .S(_04393_),
    .X(_04397_));
 sky130_fd_sc_hd__o21ai_1 _10093_ (.A1(_04181_),
    .A2(_04397_),
    .B1(_00227_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ));
 sky130_fd_sc_hd__a41o_2 _10094_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .A2(_04345_),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .A4(_04372_),
    .B1(_00249_),
    .X(_04398_));
 sky130_fd_sc_hd__mux2_1 _10095_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .A1(_00235_),
    .S(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_1 _10096_ (.A(_04399_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ));
 sky130_fd_sc_hd__mux2_1 _10097_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .A1(_00292_),
    .S(_04398_),
    .X(_04400_));
 sky130_fd_sc_hd__clkbuf_1 _10098_ (.A(_04400_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ));
 sky130_fd_sc_hd__mux2_1 _10099_ (.A0(net3858),
    .A1(_00188_),
    .S(_04398_),
    .X(_04401_));
 sky130_fd_sc_hd__clkbuf_1 _10100_ (.A(_04401_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ));
 sky130_fd_sc_hd__mux2_1 _10101_ (.A0(net4093),
    .A1(_00527_),
    .S(_04398_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _10102_ (.A(_04402_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ));
 sky130_fd_sc_hd__inv_2 _10103_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .Y(_04403_));
 sky130_fd_sc_hd__o31a_2 _10104_ (.A1(_04403_),
    .A2(_04336_),
    .A3(_04337_),
    .B1(_01497_),
    .X(_04404_));
 sky130_fd_sc_hd__mux2_1 _10105_ (.A0(_00172_),
    .A1(net4004),
    .S(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _10106_ (.A(_04405_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ));
 sky130_fd_sc_hd__mux2_1 _10107_ (.A0(_00185_),
    .A1(net3412),
    .S(_04404_),
    .X(_04406_));
 sky130_fd_sc_hd__clkbuf_1 _10108_ (.A(_04406_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ));
 sky130_fd_sc_hd__mux2_1 _10109_ (.A0(_00189_),
    .A1(net3783),
    .S(_04404_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_1 _10110_ (.A(_04407_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ));
 sky130_fd_sc_hd__mux2_1 _10111_ (.A0(_00192_),
    .A1(net3893),
    .S(_04404_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_1 _10112_ (.A(_04408_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ));
 sky130_fd_sc_hd__or2_1 _10113_ (.A(_04336_),
    .B(_04357_),
    .X(_04409_));
 sky130_fd_sc_hd__o21a_2 _10114_ (.A1(_04346_),
    .A2(_04409_),
    .B1(_01489_),
    .X(_04410_));
 sky130_fd_sc_hd__mux2_1 _10115_ (.A0(_00172_),
    .A1(net3729),
    .S(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_1 _10116_ (.A(_04411_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ));
 sky130_fd_sc_hd__mux2_1 _10117_ (.A0(_00185_),
    .A1(net3438),
    .S(_04410_),
    .X(_04412_));
 sky130_fd_sc_hd__clkbuf_1 _10118_ (.A(_04412_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ));
 sky130_fd_sc_hd__mux2_1 _10119_ (.A0(_00189_),
    .A1(net3776),
    .S(_04410_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_1 _10120_ (.A(_04413_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ));
 sky130_fd_sc_hd__mux2_1 _10121_ (.A0(_00192_),
    .A1(net3589),
    .S(_04410_),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_1 _10122_ (.A(_04414_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ));
 sky130_fd_sc_hd__nor2_2 _10123_ (.A(_04353_),
    .B(_04409_),
    .Y(_04415_));
 sky130_fd_sc_hd__mux2_1 _10124_ (.A0(_03447_),
    .A1(_04359_),
    .S(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__o21ai_1 _10125_ (.A1(_04181_),
    .A2(_04416_),
    .B1(_00237_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ));
 sky130_fd_sc_hd__buf_8 _10126_ (.A(_02637_),
    .X(_04417_));
 sky130_fd_sc_hd__mux2_1 _10127_ (.A0(_03442_),
    .A1(_04363_),
    .S(_04415_),
    .X(_04418_));
 sky130_fd_sc_hd__o21ai_1 _10128_ (.A1(_04417_),
    .A2(_04418_),
    .B1(_00305_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ));
 sky130_fd_sc_hd__buf_6 _10129_ (.A(_00195_),
    .X(_04419_));
 sky130_fd_sc_hd__nand2_1 _10130_ (.A(_04366_),
    .B(_04415_),
    .Y(_04420_));
 sky130_fd_sc_hd__or2_1 _10131_ (.A(net3312),
    .B(_04415_),
    .X(_04421_));
 sky130_fd_sc_hd__a31o_1 _10132_ (.A1(_04419_),
    .A2(_04420_),
    .A3(_04421_),
    .B1(_01851_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ));
 sky130_fd_sc_hd__nor2_1 _10133_ (.A(net4053),
    .B(_04415_),
    .Y(_04422_));
 sky130_fd_sc_hd__a211o_1 _10134_ (.A1(_04369_),
    .A2(_04415_),
    .B1(_04422_),
    .C1(_00228_),
    .X(_04423_));
 sky130_fd_sc_hd__nand2_1 _10135_ (.A(_00276_),
    .B(_04423_),
    .Y(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ));
 sky130_fd_sc_hd__and3_2 _10136_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(_04355_),
    .C(_04373_),
    .X(_04424_));
 sky130_fd_sc_hd__nor2_1 _10137_ (.A(_01971_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__a221o_1 _10138_ (.A1(_00288_),
    .A2(_04424_),
    .B1(_04425_),
    .B2(net3196),
    .C1(_00209_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ));
 sky130_fd_sc_hd__a221o_1 _10139_ (.A1(_00293_),
    .A2(_04424_),
    .B1(_04425_),
    .B2(net3146),
    .C1(_02872_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ));
 sky130_fd_sc_hd__a221o_1 _10140_ (.A1(_00295_),
    .A2(_04424_),
    .B1(_04425_),
    .B2(net3153),
    .C1(_00221_),
    .X(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ));
 sky130_fd_sc_hd__mux2_1 _10141_ (.A0(_03532_),
    .A1(_03533_),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[28] ),
    .X(_04426_));
 sky130_fd_sc_hd__inv_2 _10142_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[28] ),
    .Y(_04427_));
 sky130_fd_sc_hd__a211o_1 _10143_ (.A1(_00893_),
    .A2(_00968_),
    .B1(_04427_),
    .C1(_00971_),
    .X(_04428_));
 sky130_fd_sc_hd__inv_2 _10144_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[29] ),
    .Y(_04429_));
 sky130_fd_sc_hd__o211a_1 _10145_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[28] ),
    .A2(_03530_),
    .B1(_04428_),
    .C1(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__inv_2 _10146_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[30] ),
    .Y(_04431_));
 sky130_fd_sc_hd__a211o_1 _10147_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[29] ),
    .A2(_04426_),
    .B1(_04430_),
    .C1(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__mux4_1 _10148_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04217_),
    .A3(_04218_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[28] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[29] ),
    .X(_04433_));
 sky130_fd_sc_hd__o21a_1 _10149_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[30] ),
    .A2(_04433_),
    .B1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[31] ),
    .X(_04434_));
 sky130_fd_sc_hd__mux4_1 _10150_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[29] ),
    .S1(_04427_),
    .X(_04435_));
 sky130_fd_sc_hd__mux4_1 _10151_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[28] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[29] ),
    .X(_04436_));
 sky130_fd_sc_hd__mux2_1 _10152_ (.A0(_04435_),
    .A1(_04436_),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[30] ),
    .X(_04437_));
 sky130_fd_sc_hd__o2bb2a_1 _10153_ (.A1_N(_04432_),
    .A2_N(_04434_),
    .B1(_04437_),
    .B2(net3646),
    .X(\c.genblk1.genblk1.subs.sw.up.x.o_[7] ));
 sky130_fd_sc_hd__mux4_1 _10154_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ),
    .X(_04438_));
 sky130_fd_sc_hd__or2_1 _10155_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[26] ),
    .B(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__mux2_1 _10156_ (.A0(_03786_),
    .A1(_03787_),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ),
    .X(_04440_));
 sky130_fd_sc_hd__inv_2 _10157_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ),
    .Y(_04441_));
 sky130_fd_sc_hd__a211o_1 _10158_ (.A1(_00893_),
    .A2(_00968_),
    .B1(_04441_),
    .C1(_00971_),
    .X(_04442_));
 sky130_fd_sc_hd__inv_2 _10159_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ),
    .Y(_04443_));
 sky130_fd_sc_hd__o211a_1 _10160_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ),
    .A2(_03697_),
    .B1(_04442_),
    .C1(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__inv_2 _10161_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[26] ),
    .Y(_04445_));
 sky130_fd_sc_hd__a211o_1 _10162_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ),
    .A2(_04440_),
    .B1(_04444_),
    .C1(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__mux4_1 _10163_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ),
    .S1(_04441_),
    .X(_04447_));
 sky130_fd_sc_hd__nand2_1 _10164_ (.A(_04445_),
    .B(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__mux4_1 _10165_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ),
    .X(_04449_));
 sky130_fd_sc_hd__a21oi_1 _10166_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[26] ),
    .A2(_04449_),
    .B1(net3169),
    .Y(_04450_));
 sky130_fd_sc_hd__a32oi_1 _10167_ (.A1(net3169),
    .A2(_04439_),
    .A3(_04446_),
    .B1(_04448_),
    .B2(_04450_),
    .Y(\c.genblk1.genblk1.subs.sw.up.x.o_[6] ));
 sky130_fd_sc_hd__mux4_1 _10168_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[21] ),
    .X(_04451_));
 sky130_fd_sc_hd__or2_1 _10169_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[22] ),
    .B(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__inv_2 _10170_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[20] ),
    .Y(_04453_));
 sky130_fd_sc_hd__nand2_1 _10171_ (.A(_04453_),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .Y(_04454_));
 sky130_fd_sc_hd__a21oi_1 _10172_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[20] ),
    .A2(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .B1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[21] ),
    .Y(_04455_));
 sky130_fd_sc_hd__mux2_1 _10173_ (.A0(_03786_),
    .A1(_03787_),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[20] ),
    .X(_04456_));
 sky130_fd_sc_hd__inv_2 _10174_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[22] ),
    .Y(_04457_));
 sky130_fd_sc_hd__a221o_1 _10175_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04456_),
    .B2(\c.genblk1.genblk1.subs.sw.up.x.selects.o[21] ),
    .C1(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__mux4_1 _10176_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[21] ),
    .S1(_04453_),
    .X(_04459_));
 sky130_fd_sc_hd__nand2_1 _10177_ (.A(_04457_),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__mux4_1 _10178_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[20] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[21] ),
    .X(_04461_));
 sky130_fd_sc_hd__a21oi_1 _10179_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[22] ),
    .A2(_04461_),
    .B1(net247),
    .Y(_04462_));
 sky130_fd_sc_hd__a32oi_1 _10180_ (.A1(net247),
    .A2(_04452_),
    .A3(_04458_),
    .B1(_04460_),
    .B2(_04462_),
    .Y(\c.genblk1.genblk1.subs.sw.up.x.o_[5] ));
 sky130_fd_sc_hd__mux2_1 _10181_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[16] ),
    .X(_04463_));
 sky130_fd_sc_hd__nor2_1 _10182_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[16] ),
    .B(_03532_),
    .Y(_04464_));
 sky130_fd_sc_hd__inv_2 _10183_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[16] ),
    .Y(_04465_));
 sky130_fd_sc_hd__o21ai_1 _10184_ (.A1(_04465_),
    .A2(_03533_),
    .B1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[17] ),
    .Y(_04466_));
 sky130_fd_sc_hd__o221a_1 _10185_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[17] ),
    .A2(_04463_),
    .B1(_04464_),
    .B2(_04466_),
    .C1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[18] ),
    .X(_04467_));
 sky130_fd_sc_hd__mux4_1 _10186_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04217_),
    .A3(_04218_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[16] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[17] ),
    .X(_04468_));
 sky130_fd_sc_hd__o21ai_1 _10187_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[18] ),
    .A2(_04468_),
    .B1(net3191),
    .Y(_04469_));
 sky130_fd_sc_hd__mux4_1 _10188_ (.A0(_03780_),
    .A1(_03781_),
    .A2(_03782_),
    .A3(_03783_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[17] ),
    .S1(_04465_),
    .X(_04470_));
 sky130_fd_sc_hd__mux4_1 _10189_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[16] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[17] ),
    .X(_04471_));
 sky130_fd_sc_hd__mux2_1 _10190_ (.A0(_04470_),
    .A1(_04471_),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[18] ),
    .X(_04472_));
 sky130_fd_sc_hd__o22a_1 _10191_ (.A1(_04467_),
    .A2(_04469_),
    .B1(_04472_),
    .B2(net3191),
    .X(\c.genblk1.genblk1.subs.sw.up.x.o_[4] ));
 sky130_fd_sc_hd__nor2_1 _10192_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ),
    .B(_03532_),
    .Y(_04473_));
 sky130_fd_sc_hd__inv_2 _10193_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ),
    .Y(_04474_));
 sky130_fd_sc_hd__o21ai_1 _10194_ (.A1(_04474_),
    .A2(_03533_),
    .B1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ),
    .Y(_04475_));
 sky130_fd_sc_hd__mux2_1 _10195_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ),
    .X(_04476_));
 sky130_fd_sc_hd__o221a_1 _10196_ (.A1(_04473_),
    .A2(_04475_),
    .B1(_04476_),
    .B2(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ),
    .C1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[14] ),
    .X(_04477_));
 sky130_fd_sc_hd__mux4_1 _10197_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04217_),
    .A3(_04218_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ),
    .X(_04478_));
 sky130_fd_sc_hd__o21ai_1 _10198_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[14] ),
    .A2(_04478_),
    .B1(net3354),
    .Y(_04479_));
 sky130_fd_sc_hd__mux4_1 _10199_ (.A0(_03780_),
    .A1(_03781_),
    .A2(_03782_),
    .A3(_03783_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ),
    .S1(_04474_),
    .X(_04480_));
 sky130_fd_sc_hd__mux4_1 _10200_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ),
    .X(_04481_));
 sky130_fd_sc_hd__mux2_1 _10201_ (.A0(_04480_),
    .A1(_04481_),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[14] ),
    .X(_04482_));
 sky130_fd_sc_hd__o22a_1 _10202_ (.A1(_04477_),
    .A2(_04479_),
    .B1(_04482_),
    .B2(net3354),
    .X(\c.genblk1.genblk1.subs.sw.up.x.o_[3] ));
 sky130_fd_sc_hd__nor2_1 _10203_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ),
    .B(_03532_),
    .Y(_04483_));
 sky130_fd_sc_hd__inv_2 _10204_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ),
    .Y(_04484_));
 sky130_fd_sc_hd__o21ai_1 _10205_ (.A1(_04484_),
    .A2(_03533_),
    .B1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[9] ),
    .Y(_04485_));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ),
    .X(_04486_));
 sky130_fd_sc_hd__o221ai_1 _10207_ (.A1(_04483_),
    .A2(_04485_),
    .B1(_04486_),
    .B2(\c.genblk1.genblk1.subs.sw.up.x.selects.o[9] ),
    .C1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[10] ),
    .Y(_04487_));
 sky130_fd_sc_hd__mux4_1 _10208_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04217_),
    .A3(_04218_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[9] ),
    .X(_04488_));
 sky130_fd_sc_hd__o21a_1 _10209_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[10] ),
    .A2(_04488_),
    .B1(net3388),
    .X(_04489_));
 sky130_fd_sc_hd__mux4_1 _10210_ (.A0(_03780_),
    .A1(_03781_),
    .A2(_03782_),
    .A3(_03783_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[9] ),
    .S1(_04484_),
    .X(_04490_));
 sky130_fd_sc_hd__mux4_1 _10211_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[9] ),
    .X(_04491_));
 sky130_fd_sc_hd__mux2_1 _10212_ (.A0(_04490_),
    .A1(_04491_),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[10] ),
    .X(_04492_));
 sky130_fd_sc_hd__o2bb2a_1 _10213_ (.A1_N(_04487_),
    .A2_N(_04489_),
    .B1(_04492_),
    .B2(net3388),
    .X(\c.genblk1.genblk1.subs.sw.up.x.o_[2] ));
 sky130_fd_sc_hd__mux4_1 _10214_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ),
    .X(_04493_));
 sky130_fd_sc_hd__or2_1 _10215_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[6] ),
    .B(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__inv_2 _10216_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ),
    .Y(_04495_));
 sky130_fd_sc_hd__mux2_1 _10217_ (.A0(_03697_),
    .A1(_03698_),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ),
    .X(_04496_));
 sky130_fd_sc_hd__or2_1 _10218_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ),
    .B(_03786_),
    .X(_04497_));
 sky130_fd_sc_hd__inv_2 _10219_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ),
    .Y(_04498_));
 sky130_fd_sc_hd__o21a_1 _10220_ (.A1(_04498_),
    .A2(_03787_),
    .B1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ),
    .X(_04499_));
 sky130_fd_sc_hd__inv_2 _10221_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[6] ),
    .Y(_04500_));
 sky130_fd_sc_hd__a221o_1 _10222_ (.A1(_04495_),
    .A2(_04496_),
    .B1(_04497_),
    .B2(_04499_),
    .C1(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__mux4_1 _10223_ (.A0(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ),
    .S1(_04498_),
    .X(_04502_));
 sky130_fd_sc_hd__nand2_1 _10224_ (.A(_04500_),
    .B(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__mux4_1 _10225_ (.A0(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .A2(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .A3(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ),
    .X(_04504_));
 sky130_fd_sc_hd__a21oi_1 _10226_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[6] ),
    .A2(_04504_),
    .B1(net3215),
    .Y(_04505_));
 sky130_fd_sc_hd__a32oi_1 _10227_ (.A1(net3215),
    .A2(_04494_),
    .A3(_04501_),
    .B1(_04503_),
    .B2(_04505_),
    .Y(\c.genblk1.genblk1.subs.sw.up.x.o_[1] ));
 sky130_fd_sc_hd__nor2_1 _10228_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[0] ),
    .B(_03532_),
    .Y(_04506_));
 sky130_fd_sc_hd__inv_2 _10229_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[0] ),
    .Y(_04507_));
 sky130_fd_sc_hd__o21ai_1 _10230_ (.A1(_04507_),
    .A2(_03533_),
    .B1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[1] ),
    .Y(_04508_));
 sky130_fd_sc_hd__mux2_1 _10231_ (.A0(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .A1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[0] ),
    .X(_04509_));
 sky130_fd_sc_hd__o221a_1 _10232_ (.A1(_04506_),
    .A2(_04508_),
    .B1(_04509_),
    .B2(\c.genblk1.genblk1.subs.sw.up.x.selects.o[1] ),
    .C1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[2] ),
    .X(_04510_));
 sky130_fd_sc_hd__mux4_1 _10233_ (.A0(_04215_),
    .A1(_04216_),
    .A2(_04217_),
    .A3(_04218_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[1] ),
    .X(_04511_));
 sky130_fd_sc_hd__o21ai_1 _10234_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[2] ),
    .A2(_04511_),
    .B1(net3225),
    .Y(_04512_));
 sky130_fd_sc_hd__mux4_1 _10235_ (.A0(_03780_),
    .A1(_03781_),
    .A2(_03782_),
    .A3(_03783_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[1] ),
    .S1(_04507_),
    .X(_04513_));
 sky130_fd_sc_hd__mux4_1 _10236_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\c.genblk1.genblk1.subs.sw.up.x.selects.o[0] ),
    .S1(\c.genblk1.genblk1.subs.sw.up.x.selects.o[1] ),
    .X(_04514_));
 sky130_fd_sc_hd__mux2_1 _10237_ (.A0(_04513_),
    .A1(_04514_),
    .S(\c.genblk1.genblk1.subs.sw.up.x.selects.o[2] ),
    .X(_04515_));
 sky130_fd_sc_hd__o22a_1 _10238_ (.A1(_04510_),
    .A2(_04512_),
    .B1(_04515_),
    .B2(net3225),
    .X(\c.genblk1.genblk1.subs.sw.up.x.o_[0] ));
 sky130_fd_sc_hd__mux2_1 _10239_ (.A0(_03749_),
    .A1(_04209_),
    .S(_02524_),
    .X(_04516_));
 sky130_fd_sc_hd__clkbuf_1 _10240_ (.A(_04516_),
    .X(_00003_));
 sky130_fd_sc_hd__and3_1 _10241_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[5] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[1] ),
    .C(_00199_),
    .X(_04517_));
 sky130_fd_sc_hd__a31o_1 _10242_ (.A1(net3180),
    .A2(_00174_),
    .A3(_04517_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[0].x.cfgd ),
    .X(_04518_));
 sky130_fd_sc_hd__and2_1 _10243_ (.A(_04419_),
    .B(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__clkbuf_1 _10244_ (.A(_04519_),
    .X(_00016_));
 sky130_fd_sc_hd__buf_4 _10245_ (.A(_00236_),
    .X(_04520_));
 sky130_fd_sc_hd__and3b_1 _10246_ (.A_N(_04517_),
    .B(_00174_),
    .C(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[0] ),
    .X(_04521_));
 sky130_fd_sc_hd__nor2_1 _10247_ (.A(_04520_),
    .B(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__o21a_1 _10248_ (.A1(net3180),
    .A2(_00174_),
    .B1(_04522_),
    .X(_00017_));
 sky130_fd_sc_hd__and2_1 _10249_ (.A(net3335),
    .B(_04521_),
    .X(_04523_));
 sky130_fd_sc_hd__nor2_1 _10250_ (.A(net3335),
    .B(_04521_),
    .Y(_04524_));
 sky130_fd_sc_hd__nor3_1 _10251_ (.A(_04417_),
    .B(_04523_),
    .C(_04524_),
    .Y(_00018_));
 sky130_fd_sc_hd__and3_1 _10252_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ),
    .B(net4151),
    .C(_04521_),
    .X(_04525_));
 sky130_fd_sc_hd__nor2_1 _10253_ (.A(_04520_),
    .B(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__o21a_1 _10254_ (.A1(net3907),
    .A2(_04523_),
    .B1(_04526_),
    .X(_00019_));
 sky130_fd_sc_hd__and2_1 _10255_ (.A(_00198_),
    .B(_04525_),
    .X(_04527_));
 sky130_fd_sc_hd__nor2_1 _10256_ (.A(_04520_),
    .B(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__o21a_1 _10257_ (.A1(_00198_),
    .A2(_04525_),
    .B1(_04528_),
    .X(_00020_));
 sky130_fd_sc_hd__and3_1 _10258_ (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ),
    .B(_00198_),
    .C(_04525_),
    .X(_04529_));
 sky130_fd_sc_hd__nor2_1 _10259_ (.A(_04520_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__o21a_1 _10260_ (.A1(net3832),
    .A2(_04527_),
    .B1(_04530_),
    .X(_00021_));
 sky130_fd_sc_hd__buf_6 _10261_ (.A(_02637_),
    .X(_04531_));
 sky130_fd_sc_hd__a21oi_1 _10262_ (.A1(net3661),
    .A2(_04529_),
    .B1(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__o21a_1 _10263_ (.A1(net3661),
    .A2(_04529_),
    .B1(_04532_),
    .X(_00022_));
 sky130_fd_sc_hd__and3_1 _10264_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[5] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[1] ),
    .C(_00330_),
    .X(_04533_));
 sky130_fd_sc_hd__a31o_1 _10265_ (.A1(net4222),
    .A2(_00313_),
    .A3(_04533_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[1].x.cfgd ),
    .X(_04534_));
 sky130_fd_sc_hd__and2_1 _10266_ (.A(_04419_),
    .B(_04534_),
    .X(_04535_));
 sky130_fd_sc_hd__clkbuf_1 _10267_ (.A(_04535_),
    .X(_00023_));
 sky130_fd_sc_hd__and3b_1 _10268_ (.A_N(_04533_),
    .B(_00313_),
    .C(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[0] ),
    .X(_04536_));
 sky130_fd_sc_hd__nor2_1 _10269_ (.A(_04520_),
    .B(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__o21a_1 _10270_ (.A1(net3257),
    .A2(_00313_),
    .B1(_04537_),
    .X(_00024_));
 sky130_fd_sc_hd__and2_1 _10271_ (.A(net3377),
    .B(_04536_),
    .X(_04538_));
 sky130_fd_sc_hd__a21oi_1 _10272_ (.A1(net3257),
    .A2(_00313_),
    .B1(net3377),
    .Y(_04539_));
 sky130_fd_sc_hd__nor3_1 _10273_ (.A(_04417_),
    .B(_04538_),
    .C(_04539_),
    .Y(_00025_));
 sky130_fd_sc_hd__and3_1 _10274_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ),
    .B(net3377),
    .C(_04536_),
    .X(_04540_));
 sky130_fd_sc_hd__nor2_1 _10275_ (.A(_04520_),
    .B(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__o21a_1 _10276_ (.A1(net3824),
    .A2(_04538_),
    .B1(_04541_),
    .X(_00026_));
 sky130_fd_sc_hd__and2_1 _10277_ (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ),
    .B(_04540_),
    .X(_04542_));
 sky130_fd_sc_hd__nor2_1 _10278_ (.A(_04520_),
    .B(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__o21a_1 _10279_ (.A1(net3837),
    .A2(_04540_),
    .B1(_04543_),
    .X(_00027_));
 sky130_fd_sc_hd__and3_1 _10280_ (.A(net3566),
    .B(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ),
    .C(_04540_),
    .X(_04544_));
 sky130_fd_sc_hd__nor2_1 _10281_ (.A(_04520_),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__o21a_1 _10282_ (.A1(net3566),
    .A2(_04542_),
    .B1(_04545_),
    .X(_00028_));
 sky130_fd_sc_hd__a21oi_1 _10283_ (.A1(net3777),
    .A2(_04544_),
    .B1(_04531_),
    .Y(_04546_));
 sky130_fd_sc_hd__o21a_1 _10284_ (.A1(net3777),
    .A2(_04544_),
    .B1(_04546_),
    .X(_00029_));
 sky130_fd_sc_hd__and3_1 _10285_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[5] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[1] ),
    .C(_00444_),
    .X(_04547_));
 sky130_fd_sc_hd__a31o_1 _10286_ (.A1(net3184),
    .A2(_00427_),
    .A3(_04547_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[2].x.cfgd ),
    .X(_04548_));
 sky130_fd_sc_hd__and2_1 _10287_ (.A(_04419_),
    .B(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__clkbuf_1 _10288_ (.A(_04549_),
    .X(_00030_));
 sky130_fd_sc_hd__and3b_1 _10289_ (.A_N(_04547_),
    .B(_00427_),
    .C(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[0] ),
    .X(_04550_));
 sky130_fd_sc_hd__nor2_1 _10290_ (.A(_04520_),
    .B(_04550_),
    .Y(_04551_));
 sky130_fd_sc_hd__o21a_1 _10291_ (.A1(net3184),
    .A2(_00427_),
    .B1(_04551_),
    .X(_00031_));
 sky130_fd_sc_hd__and2_1 _10292_ (.A(net3247),
    .B(_04550_),
    .X(_04552_));
 sky130_fd_sc_hd__nor2_1 _10293_ (.A(net3247),
    .B(_04550_),
    .Y(_04553_));
 sky130_fd_sc_hd__nor3_1 _10294_ (.A(_04417_),
    .B(_04552_),
    .C(net3248),
    .Y(_00032_));
 sky130_fd_sc_hd__buf_4 _10295_ (.A(_00236_),
    .X(_04554_));
 sky130_fd_sc_hd__and3_1 _10296_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ),
    .B(net3900),
    .C(_04550_),
    .X(_04555_));
 sky130_fd_sc_hd__nor2_1 _10297_ (.A(_04554_),
    .B(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__o21a_1 _10298_ (.A1(net3746),
    .A2(_04552_),
    .B1(_04556_),
    .X(_00033_));
 sky130_fd_sc_hd__and2_1 _10299_ (.A(_00438_),
    .B(_04555_),
    .X(_04557_));
 sky130_fd_sc_hd__nor2_1 _10300_ (.A(_04554_),
    .B(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__o21a_1 _10301_ (.A1(_00438_),
    .A2(_04555_),
    .B1(_04558_),
    .X(_00034_));
 sky130_fd_sc_hd__and3_1 _10302_ (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ),
    .B(_00438_),
    .C(_04555_),
    .X(_04559_));
 sky130_fd_sc_hd__nor2_1 _10303_ (.A(_04554_),
    .B(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__o21a_1 _10304_ (.A1(net3877),
    .A2(_04557_),
    .B1(_04560_),
    .X(_00035_));
 sky130_fd_sc_hd__a21oi_1 _10305_ (.A1(net3565),
    .A2(_04559_),
    .B1(_04531_),
    .Y(_04561_));
 sky130_fd_sc_hd__o21a_1 _10306_ (.A1(net3565),
    .A2(_04559_),
    .B1(_04561_),
    .X(_00036_));
 sky130_fd_sc_hd__and3_1 _10307_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[5] ),
    .B(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[1] ),
    .C(_00563_),
    .X(_04562_));
 sky130_fd_sc_hd__a31o_1 _10308_ (.A1(net4216),
    .A2(_00542_),
    .A3(_04562_),
    .B1(\c.genblk1.genblk1.subs.sw.dns[3].x.cfgd ),
    .X(_04563_));
 sky130_fd_sc_hd__and2_1 _10309_ (.A(_04419_),
    .B(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__clkbuf_1 _10310_ (.A(_04564_),
    .X(_00037_));
 sky130_fd_sc_hd__and3b_1 _10311_ (.A_N(_04562_),
    .B(_00542_),
    .C(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[0] ),
    .X(_04565_));
 sky130_fd_sc_hd__nor2_1 _10312_ (.A(_04554_),
    .B(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__o21a_1 _10313_ (.A1(net3294),
    .A2(_00542_),
    .B1(_04566_),
    .X(_00038_));
 sky130_fd_sc_hd__and2_1 _10314_ (.A(net3367),
    .B(_04565_),
    .X(_04567_));
 sky130_fd_sc_hd__a21oi_1 _10315_ (.A1(net3294),
    .A2(_00542_),
    .B1(net3367),
    .Y(_04568_));
 sky130_fd_sc_hd__nor3_1 _10316_ (.A(_04417_),
    .B(_04567_),
    .C(_04568_),
    .Y(_00039_));
 sky130_fd_sc_hd__and3_1 _10317_ (.A(_00556_),
    .B(net4223),
    .C(_04565_),
    .X(_04569_));
 sky130_fd_sc_hd__nor2_1 _10318_ (.A(_04554_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__o21a_1 _10319_ (.A1(_00556_),
    .A2(_04567_),
    .B1(_04570_),
    .X(_00040_));
 sky130_fd_sc_hd__and2_1 _10320_ (.A(_00555_),
    .B(_04569_),
    .X(_04571_));
 sky130_fd_sc_hd__nor2_1 _10321_ (.A(_04554_),
    .B(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__o21a_1 _10322_ (.A1(_00555_),
    .A2(_04569_),
    .B1(_04572_),
    .X(_00041_));
 sky130_fd_sc_hd__and3_1 _10323_ (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ),
    .B(_00555_),
    .C(_04569_),
    .X(_04573_));
 sky130_fd_sc_hd__nor2_1 _10324_ (.A(_04554_),
    .B(_04573_),
    .Y(_04574_));
 sky130_fd_sc_hd__o21a_1 _10325_ (.A1(net3761),
    .A2(_04571_),
    .B1(_04574_),
    .X(_00042_));
 sky130_fd_sc_hd__a21oi_1 _10326_ (.A1(net3573),
    .A2(_04573_),
    .B1(_04531_),
    .Y(_04575_));
 sky130_fd_sc_hd__o21a_1 _10327_ (.A1(net3573),
    .A2(_04573_),
    .B1(_04575_),
    .X(_00043_));
 sky130_fd_sc_hd__and4_1 _10328_ (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[4] ),
    .B(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ),
    .C(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[2] ),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[1] ),
    .X(_04576_));
 sky130_fd_sc_hd__a31o_1 _10329_ (.A1(net3255),
    .A2(_00660_),
    .A3(_04576_),
    .B1(net27),
    .X(_04577_));
 sky130_fd_sc_hd__and2_1 _10330_ (.A(_04419_),
    .B(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__clkbuf_1 _10331_ (.A(_04578_),
    .X(_00044_));
 sky130_fd_sc_hd__and3b_1 _10332_ (.A_N(_04576_),
    .B(_00660_),
    .C(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[0] ),
    .X(_04579_));
 sky130_fd_sc_hd__nor2_1 _10333_ (.A(_04554_),
    .B(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__o21a_1 _10334_ (.A1(net3199),
    .A2(_00660_),
    .B1(_04580_),
    .X(_00045_));
 sky130_fd_sc_hd__and2_1 _10335_ (.A(net3795),
    .B(_04579_),
    .X(_04581_));
 sky130_fd_sc_hd__a21oi_1 _10336_ (.A1(net3199),
    .A2(_00660_),
    .B1(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[1] ),
    .Y(_04582_));
 sky130_fd_sc_hd__nor3_1 _10337_ (.A(_04417_),
    .B(_04581_),
    .C(net3200),
    .Y(_00046_));
 sky130_fd_sc_hd__and3_1 _10338_ (.A(net3765),
    .B(net3795),
    .C(_04579_),
    .X(_04583_));
 sky130_fd_sc_hd__nor2_1 _10339_ (.A(_04554_),
    .B(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__o21a_1 _10340_ (.A1(net3765),
    .A2(_04581_),
    .B1(_04584_),
    .X(_00047_));
 sky130_fd_sc_hd__buf_6 _10341_ (.A(_02637_),
    .X(_04585_));
 sky130_fd_sc_hd__a21oi_1 _10342_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ),
    .A2(_04583_),
    .B1(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__o21a_1 _10343_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ),
    .A2(_04583_),
    .B1(_04586_),
    .X(_00048_));
 sky130_fd_sc_hd__a21oi_1 _10344_ (.A1(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ),
    .A2(_04583_),
    .B1(net3041),
    .Y(_04587_));
 sky130_fd_sc_hd__nor2_1 _10345_ (.A(_00229_),
    .B(_04587_),
    .Y(_00049_));
 sky130_fd_sc_hd__or3_1 _10346_ (.A(_02759_),
    .B(_00888_),
    .C(_03993_),
    .X(_04588_));
 sky130_fd_sc_hd__o21a_1 _10347_ (.A1(net3820),
    .A2(_02525_),
    .B1(_04588_),
    .X(_00050_));
 sky130_fd_sc_hd__and3_1 _10348_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .C(_01456_),
    .X(_04589_));
 sky130_fd_sc_hd__a31o_1 _10349_ (.A1(net3177),
    .A2(_01434_),
    .A3(_04589_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .X(_04590_));
 sky130_fd_sc_hd__and2_1 _10350_ (.A(_04419_),
    .B(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__clkbuf_1 _10351_ (.A(_04591_),
    .X(_00051_));
 sky130_fd_sc_hd__and3b_1 _10352_ (.A_N(_04589_),
    .B(_01434_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ),
    .X(_04592_));
 sky130_fd_sc_hd__nor2_1 _10353_ (.A(_04554_),
    .B(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__o21a_1 _10354_ (.A1(net3177),
    .A2(_01434_),
    .B1(_04593_),
    .X(_00052_));
 sky130_fd_sc_hd__and2_1 _10355_ (.A(net3239),
    .B(_04592_),
    .X(_04594_));
 sky130_fd_sc_hd__nor2_1 _10356_ (.A(net3239),
    .B(_04592_),
    .Y(_04595_));
 sky130_fd_sc_hd__nor3_1 _10357_ (.A(_04417_),
    .B(_04594_),
    .C(net3240),
    .Y(_00053_));
 sky130_fd_sc_hd__buf_4 _10358_ (.A(_00236_),
    .X(_04596_));
 sky130_fd_sc_hd__and3_1 _10359_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .C(_04592_),
    .X(_04597_));
 sky130_fd_sc_hd__nor2_1 _10360_ (.A(_04596_),
    .B(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__o21a_1 _10361_ (.A1(net3649),
    .A2(_04594_),
    .B1(_04598_),
    .X(_00054_));
 sky130_fd_sc_hd__a21oi_1 _10362_ (.A1(_01425_),
    .A2(_04597_),
    .B1(_04585_),
    .Y(_04599_));
 sky130_fd_sc_hd__o21a_1 _10363_ (.A1(_01425_),
    .A2(_04597_),
    .B1(_04599_),
    .X(_00055_));
 sky130_fd_sc_hd__a21oi_1 _10364_ (.A1(_01425_),
    .A2(_04597_),
    .B1(_01426_),
    .Y(_04600_));
 sky130_fd_sc_hd__and3_1 _10365_ (.A(_01426_),
    .B(_01425_),
    .C(_04597_),
    .X(_04601_));
 sky130_fd_sc_hd__nor3_1 _10366_ (.A(_04417_),
    .B(_04600_),
    .C(_04601_),
    .Y(_00056_));
 sky130_fd_sc_hd__a21oi_1 _10367_ (.A1(net3517),
    .A2(_04601_),
    .B1(_04585_),
    .Y(_04602_));
 sky130_fd_sc_hd__o21a_1 _10368_ (.A1(net3517),
    .A2(_04601_),
    .B1(_04602_),
    .X(_00057_));
 sky130_fd_sc_hd__or3_1 _10369_ (.A(_02759_),
    .B(_01589_),
    .C(_03993_),
    .X(_04603_));
 sky130_fd_sc_hd__o21a_1 _10370_ (.A1(net3756),
    .A2(_02525_),
    .B1(_04603_),
    .X(_00058_));
 sky130_fd_sc_hd__and3_1 _10371_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .C(_01917_),
    .X(_04604_));
 sky130_fd_sc_hd__a31o_1 _10372_ (.A1(net4227),
    .A2(_01902_),
    .A3(_04604_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .X(_04605_));
 sky130_fd_sc_hd__and2_1 _10373_ (.A(_04419_),
    .B(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__clkbuf_1 _10374_ (.A(_04606_),
    .X(_00059_));
 sky130_fd_sc_hd__and3b_1 _10375_ (.A_N(_04604_),
    .B(_01902_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(_04607_));
 sky130_fd_sc_hd__nor2_1 _10376_ (.A(_04596_),
    .B(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__o21a_1 _10377_ (.A1(net3264),
    .A2(_01902_),
    .B1(_04608_),
    .X(_00060_));
 sky130_fd_sc_hd__and2_1 _10378_ (.A(net3374),
    .B(_04607_),
    .X(_04609_));
 sky130_fd_sc_hd__a21oi_1 _10379_ (.A1(net3264),
    .A2(_01902_),
    .B1(net3374),
    .Y(_04610_));
 sky130_fd_sc_hd__nor3_1 _10380_ (.A(_04417_),
    .B(_04609_),
    .C(_04610_),
    .Y(_00061_));
 sky130_fd_sc_hd__and3_1 _10381_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .C(_04607_),
    .X(_04611_));
 sky130_fd_sc_hd__nor2_1 _10382_ (.A(_04596_),
    .B(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__o21a_1 _10383_ (.A1(net3871),
    .A2(_04609_),
    .B1(_04612_),
    .X(_00062_));
 sky130_fd_sc_hd__a21oi_1 _10384_ (.A1(_01888_),
    .A2(_04611_),
    .B1(_04585_),
    .Y(_04613_));
 sky130_fd_sc_hd__o21a_1 _10385_ (.A1(_01888_),
    .A2(_04611_),
    .B1(_04613_),
    .X(_00063_));
 sky130_fd_sc_hd__a21oi_1 _10386_ (.A1(_01888_),
    .A2(_04611_),
    .B1(_01889_),
    .Y(_04614_));
 sky130_fd_sc_hd__and3_1 _10387_ (.A(_01889_),
    .B(_01888_),
    .C(_04611_),
    .X(_04615_));
 sky130_fd_sc_hd__nor3_1 _10388_ (.A(_04417_),
    .B(_04614_),
    .C(_04615_),
    .Y(_00064_));
 sky130_fd_sc_hd__a21oi_1 _10389_ (.A1(net3539),
    .A2(_04615_),
    .B1(_04585_),
    .Y(_04616_));
 sky130_fd_sc_hd__o21a_1 _10390_ (.A1(net3539),
    .A2(_04615_),
    .B1(_04616_),
    .X(_00065_));
 sky130_fd_sc_hd__and3_1 _10391_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ),
    .C(_02018_),
    .X(_04617_));
 sky130_fd_sc_hd__a31o_1 _10392_ (.A1(net3188),
    .A2(_01988_),
    .A3(_04617_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .X(_04618_));
 sky130_fd_sc_hd__and2_1 _10393_ (.A(_04419_),
    .B(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__clkbuf_1 _10394_ (.A(_04619_),
    .X(_00066_));
 sky130_fd_sc_hd__and3b_1 _10395_ (.A_N(_04617_),
    .B(_01988_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ),
    .X(_04620_));
 sky130_fd_sc_hd__nor2_1 _10396_ (.A(_04596_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__o21a_1 _10397_ (.A1(net3188),
    .A2(_01988_),
    .B1(_04621_),
    .X(_00067_));
 sky130_fd_sc_hd__clkbuf_4 _10398_ (.A(_02637_),
    .X(_04622_));
 sky130_fd_sc_hd__and2_1 _10399_ (.A(net3304),
    .B(_04620_),
    .X(_04623_));
 sky130_fd_sc_hd__nor2_1 _10400_ (.A(net3304),
    .B(_04620_),
    .Y(_04624_));
 sky130_fd_sc_hd__nor3_1 _10401_ (.A(_04622_),
    .B(_04623_),
    .C(_04624_),
    .Y(_00068_));
 sky130_fd_sc_hd__and3_1 _10402_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .B(net3304),
    .C(_04620_),
    .X(_04625_));
 sky130_fd_sc_hd__nor2_1 _10403_ (.A(_04596_),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__o21a_1 _10404_ (.A1(net3867),
    .A2(_04623_),
    .B1(_04626_),
    .X(_00069_));
 sky130_fd_sc_hd__a21oi_1 _10405_ (.A1(_01990_),
    .A2(_04625_),
    .B1(_04585_),
    .Y(_04627_));
 sky130_fd_sc_hd__o21a_1 _10406_ (.A1(_01990_),
    .A2(_04625_),
    .B1(_04627_),
    .X(_00070_));
 sky130_fd_sc_hd__a21oi_1 _10407_ (.A1(_01990_),
    .A2(_04625_),
    .B1(net3303),
    .Y(_04628_));
 sky130_fd_sc_hd__and3_1 _10408_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .B(_01990_),
    .C(_04625_),
    .X(_04629_));
 sky130_fd_sc_hd__nor3_1 _10409_ (.A(_04622_),
    .B(_04628_),
    .C(_04629_),
    .Y(_00071_));
 sky130_fd_sc_hd__a21oi_1 _10410_ (.A1(net3514),
    .A2(_04629_),
    .B1(_04585_),
    .Y(_04630_));
 sky130_fd_sc_hd__o21a_1 _10411_ (.A1(net3514),
    .A2(_04629_),
    .B1(_04630_),
    .X(_00072_));
 sky130_fd_sc_hd__and3_1 _10412_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .C(_02120_),
    .X(_04631_));
 sky130_fd_sc_hd__a31o_1 _10413_ (.A1(net3269),
    .A2(_02101_),
    .A3(_04631_),
    .B1(\c.genblk1.genblk1.subs.cs[3].c.cfgd ),
    .X(_04632_));
 sky130_fd_sc_hd__and2_1 _10414_ (.A(_04419_),
    .B(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__clkbuf_1 _10415_ (.A(_04633_),
    .X(_00073_));
 sky130_fd_sc_hd__and3b_1 _10416_ (.A_N(_04631_),
    .B(_02101_),
    .C(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(_04634_));
 sky130_fd_sc_hd__nor2_1 _10417_ (.A(_04596_),
    .B(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__o21a_1 _10418_ (.A1(net3269),
    .A2(_02101_),
    .B1(_04635_),
    .X(_00074_));
 sky130_fd_sc_hd__and2_1 _10419_ (.A(net3348),
    .B(_04634_),
    .X(_04636_));
 sky130_fd_sc_hd__a21oi_1 _10420_ (.A1(net3269),
    .A2(_02101_),
    .B1(net3348),
    .Y(_04637_));
 sky130_fd_sc_hd__nor3_1 _10421_ (.A(_04622_),
    .B(_04636_),
    .C(_04637_),
    .Y(_00075_));
 sky130_fd_sc_hd__and3_1 _10422_ (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .B(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .C(_04634_),
    .X(_04638_));
 sky130_fd_sc_hd__nor2_1 _10423_ (.A(_04596_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__o21a_1 _10424_ (.A1(net3636),
    .A2(_04636_),
    .B1(_04639_),
    .X(_00076_));
 sky130_fd_sc_hd__a21oi_1 _10425_ (.A1(_02088_),
    .A2(_04638_),
    .B1(_04585_),
    .Y(_04640_));
 sky130_fd_sc_hd__o21a_1 _10426_ (.A1(_02088_),
    .A2(_04638_),
    .B1(_04640_),
    .X(_00077_));
 sky130_fd_sc_hd__a21oi_1 _10427_ (.A1(_02088_),
    .A2(_04638_),
    .B1(_02089_),
    .Y(_04641_));
 sky130_fd_sc_hd__and3_1 _10428_ (.A(_02089_),
    .B(_02088_),
    .C(_04638_),
    .X(_04642_));
 sky130_fd_sc_hd__nor3_1 _10429_ (.A(_04622_),
    .B(_04641_),
    .C(_04642_),
    .Y(_00078_));
 sky130_fd_sc_hd__a21oi_1 _10430_ (.A1(net3533),
    .A2(_04642_),
    .B1(_04585_),
    .Y(_04643_));
 sky130_fd_sc_hd__o21a_1 _10431_ (.A1(net3533),
    .A2(_04642_),
    .B1(_04643_),
    .X(_00079_));
 sky130_fd_sc_hd__or3_1 _10432_ (.A(_02759_),
    .B(_00889_),
    .C(_03993_),
    .X(_04644_));
 sky130_fd_sc_hd__o21a_1 _10433_ (.A1(net3884),
    .A2(_02525_),
    .B1(_04644_),
    .X(_00080_));
 sky130_fd_sc_hd__buf_4 _10434_ (.A(_00195_),
    .X(_04645_));
 sky130_fd_sc_hd__and3_1 _10435_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .C(_02581_),
    .X(_04646_));
 sky130_fd_sc_hd__a31o_1 _10436_ (.A1(net3190),
    .A2(_02562_),
    .A3(_04646_),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .X(_04647_));
 sky130_fd_sc_hd__and2_1 _10437_ (.A(_04645_),
    .B(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__clkbuf_1 _10438_ (.A(_04648_),
    .X(_00081_));
 sky130_fd_sc_hd__and3b_1 _10439_ (.A_N(_04646_),
    .B(_02562_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ),
    .X(_04649_));
 sky130_fd_sc_hd__nor2_1 _10440_ (.A(_04596_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__o21a_1 _10441_ (.A1(net3190),
    .A2(_02562_),
    .B1(_04650_),
    .X(_00082_));
 sky130_fd_sc_hd__and2_1 _10442_ (.A(net3278),
    .B(_04649_),
    .X(_04651_));
 sky130_fd_sc_hd__nor2_1 _10443_ (.A(net3278),
    .B(_04649_),
    .Y(_04652_));
 sky130_fd_sc_hd__nor3_1 _10444_ (.A(_04622_),
    .B(_04651_),
    .C(net3279),
    .Y(_00083_));
 sky130_fd_sc_hd__and3_1 _10445_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .B(net3857),
    .C(_04649_),
    .X(_04653_));
 sky130_fd_sc_hd__nor2_1 _10446_ (.A(_04596_),
    .B(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__o21a_1 _10447_ (.A1(net3757),
    .A2(_04651_),
    .B1(_04654_),
    .X(_00084_));
 sky130_fd_sc_hd__a21oi_1 _10448_ (.A1(_02550_),
    .A2(_04653_),
    .B1(_04585_),
    .Y(_04655_));
 sky130_fd_sc_hd__o21a_1 _10449_ (.A1(_02550_),
    .A2(_04653_),
    .B1(_04655_),
    .X(_00085_));
 sky130_fd_sc_hd__a21oi_1 _10450_ (.A1(_02550_),
    .A2(_04653_),
    .B1(_02551_),
    .Y(_04656_));
 sky130_fd_sc_hd__and3_1 _10451_ (.A(_02551_),
    .B(_02550_),
    .C(_04653_),
    .X(_04657_));
 sky130_fd_sc_hd__nor3_1 _10452_ (.A(_04622_),
    .B(_04656_),
    .C(_04657_),
    .Y(_00086_));
 sky130_fd_sc_hd__clkbuf_8 _10453_ (.A(_00236_),
    .X(_04658_));
 sky130_fd_sc_hd__a21oi_1 _10454_ (.A1(net3784),
    .A2(_04657_),
    .B1(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__o21a_1 _10455_ (.A1(net3784),
    .A2(_04657_),
    .B1(_04659_),
    .X(_00087_));
 sky130_fd_sc_hd__or3_1 _10456_ (.A(_02759_),
    .B(_02233_),
    .C(_03993_),
    .X(_04660_));
 sky130_fd_sc_hd__o21a_1 _10457_ (.A1(net3431),
    .A2(_02525_),
    .B1(_04660_),
    .X(_00088_));
 sky130_fd_sc_hd__and3_1 _10458_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .C(_02685_),
    .X(_04661_));
 sky130_fd_sc_hd__a31o_1 _10459_ (.A1(net4228),
    .A2(_02667_),
    .A3(_04661_),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .X(_04662_));
 sky130_fd_sc_hd__and2_1 _10460_ (.A(_04645_),
    .B(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__clkbuf_1 _10461_ (.A(_04663_),
    .X(_00089_));
 sky130_fd_sc_hd__and3b_1 _10462_ (.A_N(_04661_),
    .B(_02667_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(_04664_));
 sky130_fd_sc_hd__nor2_1 _10463_ (.A(_04596_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__o21a_1 _10464_ (.A1(net3277),
    .A2(_02667_),
    .B1(_04665_),
    .X(_00090_));
 sky130_fd_sc_hd__and2_1 _10465_ (.A(net3298),
    .B(_04664_),
    .X(_04666_));
 sky130_fd_sc_hd__a21oi_1 _10466_ (.A1(net3277),
    .A2(_02667_),
    .B1(net3298),
    .Y(_04667_));
 sky130_fd_sc_hd__nor3_1 _10467_ (.A(_04622_),
    .B(_04666_),
    .C(_04667_),
    .Y(_00091_));
 sky130_fd_sc_hd__clkbuf_8 _10468_ (.A(_00236_),
    .X(_04668_));
 sky130_fd_sc_hd__and3_1 _10469_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .B(net3880),
    .C(_04664_),
    .X(_04669_));
 sky130_fd_sc_hd__nor2_1 _10470_ (.A(_04668_),
    .B(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__o21a_1 _10471_ (.A1(net3406),
    .A2(_04666_),
    .B1(_04670_),
    .X(_00092_));
 sky130_fd_sc_hd__a21oi_1 _10472_ (.A1(_02655_),
    .A2(_04669_),
    .B1(_04658_),
    .Y(_04671_));
 sky130_fd_sc_hd__o21a_1 _10473_ (.A1(_02655_),
    .A2(_04669_),
    .B1(_04671_),
    .X(_00093_));
 sky130_fd_sc_hd__a21oi_1 _10474_ (.A1(_02655_),
    .A2(_04669_),
    .B1(_02656_),
    .Y(_04672_));
 sky130_fd_sc_hd__and3_1 _10475_ (.A(_02656_),
    .B(_02655_),
    .C(_04669_),
    .X(_04673_));
 sky130_fd_sc_hd__nor3_1 _10476_ (.A(_04622_),
    .B(_04672_),
    .C(_04673_),
    .Y(_00094_));
 sky130_fd_sc_hd__a21oi_1 _10477_ (.A1(net3652),
    .A2(_04673_),
    .B1(_04658_),
    .Y(_04674_));
 sky130_fd_sc_hd__o21a_1 _10478_ (.A1(net3652),
    .A2(_04673_),
    .B1(_04674_),
    .X(_00095_));
 sky130_fd_sc_hd__and3_1 _10479_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ),
    .C(_02801_),
    .X(_04675_));
 sky130_fd_sc_hd__a31o_1 _10480_ (.A1(net4229),
    .A2(_02783_),
    .A3(_04675_),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .X(_04676_));
 sky130_fd_sc_hd__and2_1 _10481_ (.A(_04645_),
    .B(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__clkbuf_1 _10482_ (.A(_04677_),
    .X(_00096_));
 sky130_fd_sc_hd__and3b_1 _10483_ (.A_N(_04675_),
    .B(_02783_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ),
    .X(_04678_));
 sky130_fd_sc_hd__nor2_1 _10484_ (.A(_04668_),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__o21a_1 _10485_ (.A1(net3208),
    .A2(_02783_),
    .B1(_04679_),
    .X(_00097_));
 sky130_fd_sc_hd__and2_1 _10486_ (.A(net3266),
    .B(_04678_),
    .X(_04680_));
 sky130_fd_sc_hd__nor2_1 _10487_ (.A(net3266),
    .B(_04678_),
    .Y(_04681_));
 sky130_fd_sc_hd__nor3_1 _10488_ (.A(_04622_),
    .B(_04680_),
    .C(net3267),
    .Y(_00098_));
 sky130_fd_sc_hd__and3_1 _10489_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ),
    .C(_04678_),
    .X(_04682_));
 sky130_fd_sc_hd__nor2_1 _10490_ (.A(_04668_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__o21a_1 _10491_ (.A1(net3862),
    .A2(_04680_),
    .B1(_04683_),
    .X(_00099_));
 sky130_fd_sc_hd__a21oi_1 _10492_ (.A1(_02771_),
    .A2(_04682_),
    .B1(_04658_),
    .Y(_04684_));
 sky130_fd_sc_hd__o21a_1 _10493_ (.A1(_02771_),
    .A2(_04682_),
    .B1(_04684_),
    .X(_00100_));
 sky130_fd_sc_hd__a21oi_1 _10494_ (.A1(_02771_),
    .A2(_04682_),
    .B1(_02772_),
    .Y(_04685_));
 sky130_fd_sc_hd__and3_1 _10495_ (.A(_02772_),
    .B(_02771_),
    .C(_04682_),
    .X(_04686_));
 sky130_fd_sc_hd__nor3_1 _10496_ (.A(_04622_),
    .B(_04685_),
    .C(_04686_),
    .Y(_00101_));
 sky130_fd_sc_hd__a21oi_1 _10497_ (.A1(net3629),
    .A2(_04686_),
    .B1(_04658_),
    .Y(_04687_));
 sky130_fd_sc_hd__o21a_1 _10498_ (.A1(net3629),
    .A2(_04686_),
    .B1(_04687_),
    .X(_00102_));
 sky130_fd_sc_hd__and3_1 _10499_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .C(_02930_),
    .X(_04688_));
 sky130_fd_sc_hd__a31o_1 _10500_ (.A1(net4230),
    .A2(_02911_),
    .A3(_04688_),
    .B1(\c.genblk1.genblk1.subs.cs[2].c.cfgd ),
    .X(_04689_));
 sky130_fd_sc_hd__and2_1 _10501_ (.A(_04645_),
    .B(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__clkbuf_1 _10502_ (.A(_04690_),
    .X(_00103_));
 sky130_fd_sc_hd__and3b_1 _10503_ (.A_N(_04688_),
    .B(_02911_),
    .C(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(_04691_));
 sky130_fd_sc_hd__nor2_1 _10504_ (.A(_04668_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__o21a_1 _10505_ (.A1(net3251),
    .A2(_02911_),
    .B1(_04692_),
    .X(_00104_));
 sky130_fd_sc_hd__buf_4 _10506_ (.A(_02637_),
    .X(_04693_));
 sky130_fd_sc_hd__and2_1 _10507_ (.A(net3378),
    .B(_04691_),
    .X(_04694_));
 sky130_fd_sc_hd__a21oi_1 _10508_ (.A1(net3251),
    .A2(_02911_),
    .B1(net3378),
    .Y(_04695_));
 sky130_fd_sc_hd__nor3_1 _10509_ (.A(_04693_),
    .B(_04694_),
    .C(_04695_),
    .Y(_00105_));
 sky130_fd_sc_hd__and3_1 _10510_ (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .B(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .C(_04691_),
    .X(_04696_));
 sky130_fd_sc_hd__nor2_1 _10511_ (.A(_04668_),
    .B(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__o21a_1 _10512_ (.A1(net3713),
    .A2(_04694_),
    .B1(_04697_),
    .X(_00106_));
 sky130_fd_sc_hd__a21oi_1 _10513_ (.A1(_02899_),
    .A2(_04696_),
    .B1(_04658_),
    .Y(_04698_));
 sky130_fd_sc_hd__o21a_1 _10514_ (.A1(_02899_),
    .A2(_04696_),
    .B1(_04698_),
    .X(_00107_));
 sky130_fd_sc_hd__a21oi_1 _10515_ (.A1(_02899_),
    .A2(_04696_),
    .B1(_02900_),
    .Y(_04699_));
 sky130_fd_sc_hd__and3_1 _10516_ (.A(_02900_),
    .B(_02899_),
    .C(_04696_),
    .X(_04700_));
 sky130_fd_sc_hd__nor3_1 _10517_ (.A(_04693_),
    .B(_04699_),
    .C(_04700_),
    .Y(_00108_));
 sky130_fd_sc_hd__a21oi_1 _10518_ (.A1(net3443),
    .A2(_04700_),
    .B1(_04658_),
    .Y(_04701_));
 sky130_fd_sc_hd__o21a_1 _10519_ (.A1(net3443),
    .A2(_04700_),
    .B1(_04701_),
    .X(_00109_));
 sky130_fd_sc_hd__or3_1 _10520_ (.A(_02759_),
    .B(_01590_),
    .C(_03993_),
    .X(_04702_));
 sky130_fd_sc_hd__o21a_1 _10521_ (.A1(net3864),
    .A2(_02525_),
    .B1(_04702_),
    .X(_00110_));
 sky130_fd_sc_hd__and3_1 _10522_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .C(_03038_),
    .X(_04703_));
 sky130_fd_sc_hd__a31o_1 _10523_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ),
    .A2(_03022_),
    .A3(_04703_),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .X(_04704_));
 sky130_fd_sc_hd__and2_1 _10524_ (.A(_04645_),
    .B(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__clkbuf_1 _10525_ (.A(_04705_),
    .X(_00111_));
 sky130_fd_sc_hd__and3b_1 _10526_ (.A_N(_04703_),
    .B(_03022_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ),
    .X(_04706_));
 sky130_fd_sc_hd__nor2_1 _10527_ (.A(_04668_),
    .B(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__o21a_1 _10528_ (.A1(net3189),
    .A2(_03022_),
    .B1(_04707_),
    .X(_00112_));
 sky130_fd_sc_hd__and2_1 _10529_ (.A(net3252),
    .B(_04706_),
    .X(_04708_));
 sky130_fd_sc_hd__nor2_1 _10530_ (.A(net3252),
    .B(_04706_),
    .Y(_04709_));
 sky130_fd_sc_hd__nor3_1 _10531_ (.A(_04693_),
    .B(_04708_),
    .C(_04709_),
    .Y(_00113_));
 sky130_fd_sc_hd__and3_1 _10532_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .C(_04706_),
    .X(_04710_));
 sky130_fd_sc_hd__nor2_1 _10533_ (.A(_04668_),
    .B(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__o21a_1 _10534_ (.A1(net3584),
    .A2(_04708_),
    .B1(_04711_),
    .X(_00114_));
 sky130_fd_sc_hd__a21oi_1 _10535_ (.A1(_03009_),
    .A2(_04710_),
    .B1(_04658_),
    .Y(_04712_));
 sky130_fd_sc_hd__o21a_1 _10536_ (.A1(_03009_),
    .A2(_04710_),
    .B1(_04712_),
    .X(_00115_));
 sky130_fd_sc_hd__a21oi_1 _10537_ (.A1(_03009_),
    .A2(_04710_),
    .B1(_03010_),
    .Y(_04713_));
 sky130_fd_sc_hd__and3_1 _10538_ (.A(_03010_),
    .B(_03009_),
    .C(_04710_),
    .X(_04714_));
 sky130_fd_sc_hd__nor3_1 _10539_ (.A(_04693_),
    .B(_04713_),
    .C(_04714_),
    .Y(_00116_));
 sky130_fd_sc_hd__a21oi_1 _10540_ (.A1(net3473),
    .A2(_04714_),
    .B1(_04658_),
    .Y(_04715_));
 sky130_fd_sc_hd__o21a_1 _10541_ (.A1(net3473),
    .A2(_04714_),
    .B1(_04715_),
    .X(_00117_));
 sky130_fd_sc_hd__or3_1 _10542_ (.A(_02759_),
    .B(_00792_),
    .C(_03993_),
    .X(_04716_));
 sky130_fd_sc_hd__o21a_1 _10543_ (.A1(net3730),
    .A2(_02525_),
    .B1(_04716_),
    .X(_00118_));
 sky130_fd_sc_hd__and3_1 _10544_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .C(_03152_),
    .X(_04717_));
 sky130_fd_sc_hd__a31o_1 _10545_ (.A1(net4217),
    .A2(_03133_),
    .A3(_04717_),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .X(_04718_));
 sky130_fd_sc_hd__and2_1 _10546_ (.A(_04645_),
    .B(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__clkbuf_1 _10547_ (.A(_04719_),
    .X(_00119_));
 sky130_fd_sc_hd__and3b_1 _10548_ (.A_N(_04717_),
    .B(_03133_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(_04720_));
 sky130_fd_sc_hd__nor2_1 _10549_ (.A(_04668_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__o21a_1 _10550_ (.A1(net3249),
    .A2(_03133_),
    .B1(_04721_),
    .X(_00120_));
 sky130_fd_sc_hd__and2_1 _10551_ (.A(net3323),
    .B(_04720_),
    .X(_04722_));
 sky130_fd_sc_hd__a21oi_1 _10552_ (.A1(net3249),
    .A2(_03133_),
    .B1(net3323),
    .Y(_04723_));
 sky130_fd_sc_hd__nor3_1 _10553_ (.A(_04693_),
    .B(_04722_),
    .C(_04723_),
    .Y(_00121_));
 sky130_fd_sc_hd__and3_1 _10554_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .C(_04720_),
    .X(_04724_));
 sky130_fd_sc_hd__nor2_1 _10555_ (.A(_04668_),
    .B(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__o21a_1 _10556_ (.A1(net3599),
    .A2(_04722_),
    .B1(_04725_),
    .X(_00122_));
 sky130_fd_sc_hd__a21oi_1 _10557_ (.A1(_03121_),
    .A2(_04724_),
    .B1(_04658_),
    .Y(_04726_));
 sky130_fd_sc_hd__o21a_1 _10558_ (.A1(_03121_),
    .A2(_04724_),
    .B1(_04726_),
    .X(_00123_));
 sky130_fd_sc_hd__a21oi_1 _10559_ (.A1(_03121_),
    .A2(_04724_),
    .B1(_03122_),
    .Y(_04727_));
 sky130_fd_sc_hd__and3_1 _10560_ (.A(_03122_),
    .B(_03121_),
    .C(_04724_),
    .X(_04728_));
 sky130_fd_sc_hd__nor3_1 _10561_ (.A(_04693_),
    .B(_04727_),
    .C(_04728_),
    .Y(_00124_));
 sky130_fd_sc_hd__buf_6 _10562_ (.A(_00236_),
    .X(_04729_));
 sky130_fd_sc_hd__a21oi_1 _10563_ (.A1(net3550),
    .A2(_04728_),
    .B1(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__o21a_1 _10564_ (.A1(net3550),
    .A2(_04728_),
    .B1(_04730_),
    .X(_00125_));
 sky130_fd_sc_hd__and3_1 _10565_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ),
    .C(_03269_),
    .X(_04731_));
 sky130_fd_sc_hd__a31o_1 _10566_ (.A1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ),
    .A2(_03250_),
    .A3(_04731_),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .X(_04732_));
 sky130_fd_sc_hd__and2_1 _10567_ (.A(_04645_),
    .B(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__clkbuf_1 _10568_ (.A(_04733_),
    .X(_00126_));
 sky130_fd_sc_hd__and3b_1 _10569_ (.A_N(_04731_),
    .B(_03250_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ),
    .X(_04734_));
 sky130_fd_sc_hd__nor2_1 _10570_ (.A(_04668_),
    .B(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__o21a_1 _10571_ (.A1(net3193),
    .A2(_03250_),
    .B1(_04735_),
    .X(_00127_));
 sky130_fd_sc_hd__and2_1 _10572_ (.A(net3237),
    .B(_04734_),
    .X(_04736_));
 sky130_fd_sc_hd__nor2_1 _10573_ (.A(net3237),
    .B(_04734_),
    .Y(_04737_));
 sky130_fd_sc_hd__nor3_1 _10574_ (.A(_04693_),
    .B(_04736_),
    .C(_04737_),
    .Y(_00128_));
 sky130_fd_sc_hd__buf_4 _10575_ (.A(_00236_),
    .X(_04738_));
 sky130_fd_sc_hd__and3_1 _10576_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .B(net3237),
    .C(_04734_),
    .X(_04739_));
 sky130_fd_sc_hd__nor2_1 _10577_ (.A(_04738_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__o21a_1 _10578_ (.A1(net3902),
    .A2(_04736_),
    .B1(_04740_),
    .X(_00129_));
 sky130_fd_sc_hd__and2_1 _10579_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .B(_04739_),
    .X(_04741_));
 sky130_fd_sc_hd__nor2_1 _10580_ (.A(_04738_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__o21a_1 _10581_ (.A1(net3463),
    .A2(_04739_),
    .B1(_04742_),
    .X(_00130_));
 sky130_fd_sc_hd__a21oi_1 _10582_ (.A1(_03239_),
    .A2(_04741_),
    .B1(_04729_),
    .Y(_04743_));
 sky130_fd_sc_hd__o21a_1 _10583_ (.A1(_03239_),
    .A2(_04741_),
    .B1(_04743_),
    .X(_00131_));
 sky130_fd_sc_hd__a21oi_1 _10584_ (.A1(_03239_),
    .A2(_04741_),
    .B1(net3592),
    .Y(_04744_));
 sky130_fd_sc_hd__a31o_1 _10585_ (.A1(net3592),
    .A2(_03239_),
    .A3(_04741_),
    .B1(_00228_),
    .X(_04745_));
 sky130_fd_sc_hd__nor2_1 _10586_ (.A(_04744_),
    .B(_04745_),
    .Y(_00132_));
 sky130_fd_sc_hd__and3_1 _10587_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .C(_03387_),
    .X(_04746_));
 sky130_fd_sc_hd__a31o_1 _10588_ (.A1(net4220),
    .A2(_03368_),
    .A3(_04746_),
    .B1(\c.genblk1.genblk1.subs.cs[1].c.cfgd ),
    .X(_04747_));
 sky130_fd_sc_hd__and2_1 _10589_ (.A(_04645_),
    .B(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__clkbuf_1 _10590_ (.A(_04748_),
    .X(_00133_));
 sky130_fd_sc_hd__and3b_1 _10591_ (.A_N(_04746_),
    .B(_03368_),
    .C(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(_04749_));
 sky130_fd_sc_hd__nor2_1 _10592_ (.A(_04738_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__o21a_1 _10593_ (.A1(net3265),
    .A2(_03368_),
    .B1(_04750_),
    .X(_00134_));
 sky130_fd_sc_hd__and2_1 _10594_ (.A(net3371),
    .B(_04749_),
    .X(_04751_));
 sky130_fd_sc_hd__a21oi_1 _10595_ (.A1(net3265),
    .A2(_03368_),
    .B1(net3371),
    .Y(_04752_));
 sky130_fd_sc_hd__nor3_1 _10596_ (.A(_04693_),
    .B(_04751_),
    .C(_04752_),
    .Y(_00135_));
 sky130_fd_sc_hd__and3_1 _10597_ (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .B(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .C(_04749_),
    .X(_04753_));
 sky130_fd_sc_hd__nor2_1 _10598_ (.A(_04738_),
    .B(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__o21a_1 _10599_ (.A1(net3471),
    .A2(_04751_),
    .B1(_04754_),
    .X(_00136_));
 sky130_fd_sc_hd__a21oi_1 _10600_ (.A1(_03356_),
    .A2(_04753_),
    .B1(_04729_),
    .Y(_04755_));
 sky130_fd_sc_hd__o21a_1 _10601_ (.A1(_03356_),
    .A2(_04753_),
    .B1(_04755_),
    .X(_00137_));
 sky130_fd_sc_hd__a21oi_1 _10602_ (.A1(_03356_),
    .A2(_04753_),
    .B1(_03357_),
    .Y(_04756_));
 sky130_fd_sc_hd__and3_1 _10603_ (.A(_03357_),
    .B(_03356_),
    .C(_04753_),
    .X(_04757_));
 sky130_fd_sc_hd__nor3_1 _10604_ (.A(_04693_),
    .B(_04756_),
    .C(_04757_),
    .Y(_00138_));
 sky130_fd_sc_hd__a21oi_1 _10605_ (.A1(net3712),
    .A2(_04757_),
    .B1(_04729_),
    .Y(_04758_));
 sky130_fd_sc_hd__o21a_1 _10606_ (.A1(net3712),
    .A2(_04757_),
    .B1(_04758_),
    .X(_00139_));
 sky130_fd_sc_hd__or3_1 _10607_ (.A(_02759_),
    .B(_02234_),
    .C(_03993_),
    .X(_04759_));
 sky130_fd_sc_hd__o21a_1 _10608_ (.A1(net3426),
    .A2(_02525_),
    .B1(_04759_),
    .X(_00140_));
 sky130_fd_sc_hd__and3_1 _10609_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .C(_03644_),
    .X(_04760_));
 sky130_fd_sc_hd__a31o_1 _10610_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ),
    .A2(_03624_),
    .A3(_04760_),
    .B1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ),
    .X(_04761_));
 sky130_fd_sc_hd__and2_1 _10611_ (.A(_04645_),
    .B(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__clkbuf_1 _10612_ (.A(_04762_),
    .X(_00141_));
 sky130_fd_sc_hd__and3b_1 _10613_ (.A_N(_04760_),
    .B(_03624_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ),
    .X(_04763_));
 sky130_fd_sc_hd__nor2_1 _10614_ (.A(_04738_),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__o21a_1 _10615_ (.A1(net3182),
    .A2(_03624_),
    .B1(_04764_),
    .X(_00142_));
 sky130_fd_sc_hd__and2_1 _10616_ (.A(net3268),
    .B(_04763_),
    .X(_04765_));
 sky130_fd_sc_hd__nor2_1 _10617_ (.A(net3268),
    .B(_04763_),
    .Y(_04766_));
 sky130_fd_sc_hd__nor3_1 _10618_ (.A(_04693_),
    .B(_04765_),
    .C(_04766_),
    .Y(_00143_));
 sky130_fd_sc_hd__and3_1 _10619_ (.A(net3670),
    .B(net3268),
    .C(_04763_),
    .X(_04767_));
 sky130_fd_sc_hd__nor2_1 _10620_ (.A(_04738_),
    .B(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__o21a_1 _10621_ (.A1(net3670),
    .A2(_04765_),
    .B1(_04768_),
    .X(_00144_));
 sky130_fd_sc_hd__a21oi_1 _10622_ (.A1(_03614_),
    .A2(_04767_),
    .B1(_04729_),
    .Y(_04769_));
 sky130_fd_sc_hd__o21a_1 _10623_ (.A1(_03614_),
    .A2(_04767_),
    .B1(_04769_),
    .X(_00145_));
 sky130_fd_sc_hd__a21oi_1 _10624_ (.A1(_03614_),
    .A2(_04767_),
    .B1(_03615_),
    .Y(_04770_));
 sky130_fd_sc_hd__and3_1 _10625_ (.A(_03615_),
    .B(_03614_),
    .C(_04767_),
    .X(_04771_));
 sky130_fd_sc_hd__nor3_1 _10626_ (.A(_04531_),
    .B(_04770_),
    .C(_04771_),
    .Y(_00146_));
 sky130_fd_sc_hd__a21oi_1 _10627_ (.A1(net3887),
    .A2(_04771_),
    .B1(_04729_),
    .Y(_04772_));
 sky130_fd_sc_hd__o21a_1 _10628_ (.A1(net3887),
    .A2(_04771_),
    .B1(_04772_),
    .X(_00147_));
 sky130_fd_sc_hd__and3_1 _10629_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .C(_03922_),
    .X(_04773_));
 sky130_fd_sc_hd__a31o_1 _10630_ (.A1(net4221),
    .A2(_03903_),
    .A3(_04773_),
    .B1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ),
    .X(_04774_));
 sky130_fd_sc_hd__and2_1 _10631_ (.A(_04645_),
    .B(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__clkbuf_1 _10632_ (.A(_04775_),
    .X(_00148_));
 sky130_fd_sc_hd__and3b_1 _10633_ (.A_N(_04773_),
    .B(_03903_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(_04776_));
 sky130_fd_sc_hd__nor2_1 _10634_ (.A(_04738_),
    .B(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__o21a_1 _10635_ (.A1(net3280),
    .A2(_03903_),
    .B1(_04777_),
    .X(_00149_));
 sky130_fd_sc_hd__and2_1 _10636_ (.A(net3375),
    .B(_04776_),
    .X(_04778_));
 sky130_fd_sc_hd__a21oi_1 _10637_ (.A1(net3280),
    .A2(_03903_),
    .B1(net3375),
    .Y(_04779_));
 sky130_fd_sc_hd__nor3_1 _10638_ (.A(_04531_),
    .B(_04778_),
    .C(_04779_),
    .Y(_00150_));
 sky130_fd_sc_hd__and3_1 _10639_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .B(net3375),
    .C(_04776_),
    .X(_04780_));
 sky130_fd_sc_hd__nor2_1 _10640_ (.A(_04738_),
    .B(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__o21a_1 _10641_ (.A1(net3892),
    .A2(_04778_),
    .B1(_04781_),
    .X(_00151_));
 sky130_fd_sc_hd__a21oi_1 _10642_ (.A1(_03877_),
    .A2(_04780_),
    .B1(_04729_),
    .Y(_04782_));
 sky130_fd_sc_hd__o21a_1 _10643_ (.A1(_03877_),
    .A2(_04780_),
    .B1(_04782_),
    .X(_00152_));
 sky130_fd_sc_hd__a21oi_1 _10644_ (.A1(_03877_),
    .A2(_04780_),
    .B1(_03878_),
    .Y(_04783_));
 sky130_fd_sc_hd__and3_1 _10645_ (.A(_03878_),
    .B(_03877_),
    .C(_04780_),
    .X(_04784_));
 sky130_fd_sc_hd__nor3_1 _10646_ (.A(_04531_),
    .B(_04783_),
    .C(_04784_),
    .Y(_00153_));
 sky130_fd_sc_hd__a21oi_1 _10647_ (.A1(net3621),
    .A2(_04784_),
    .B1(_04729_),
    .Y(_04785_));
 sky130_fd_sc_hd__o21a_1 _10648_ (.A1(net3621),
    .A2(_04784_),
    .B1(_04785_),
    .X(_00154_));
 sky130_fd_sc_hd__and3_1 _10649_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ),
    .C(_04155_),
    .X(_04786_));
 sky130_fd_sc_hd__a31o_1 _10650_ (.A1(net3179),
    .A2(_04135_),
    .A3(_04786_),
    .B1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ),
    .X(_04787_));
 sky130_fd_sc_hd__and2_1 _10651_ (.A(_00196_),
    .B(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__clkbuf_1 _10652_ (.A(_04788_),
    .X(_00155_));
 sky130_fd_sc_hd__and3b_1 _10653_ (.A_N(_04786_),
    .B(_04135_),
    .C(net3179),
    .X(_04789_));
 sky130_fd_sc_hd__nor2_1 _10654_ (.A(_04738_),
    .B(_04789_),
    .Y(_04790_));
 sky130_fd_sc_hd__o21a_1 _10655_ (.A1(net3179),
    .A2(_04135_),
    .B1(_04790_),
    .X(_00156_));
 sky130_fd_sc_hd__and2_1 _10656_ (.A(net3261),
    .B(_04789_),
    .X(_04791_));
 sky130_fd_sc_hd__nor2_1 _10657_ (.A(net3261),
    .B(_04789_),
    .Y(_04792_));
 sky130_fd_sc_hd__nor3_1 _10658_ (.A(_04531_),
    .B(_04791_),
    .C(_04792_),
    .Y(_00157_));
 sky130_fd_sc_hd__and3_1 _10659_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ),
    .C(_04789_),
    .X(_04793_));
 sky130_fd_sc_hd__nor2_1 _10660_ (.A(_04738_),
    .B(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__o21a_1 _10661_ (.A1(net3878),
    .A2(_04791_),
    .B1(_04794_),
    .X(_00158_));
 sky130_fd_sc_hd__and2_1 _10662_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .B(_04793_),
    .X(_04795_));
 sky130_fd_sc_hd__nor2_1 _10663_ (.A(_00268_),
    .B(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__o21a_1 _10664_ (.A1(net3446),
    .A2(_04793_),
    .B1(_04796_),
    .X(_00159_));
 sky130_fd_sc_hd__a21oi_1 _10665_ (.A1(_04127_),
    .A2(_04795_),
    .B1(_04729_),
    .Y(_04797_));
 sky130_fd_sc_hd__o21a_1 _10666_ (.A1(_04127_),
    .A2(_04795_),
    .B1(_04797_),
    .X(_00160_));
 sky130_fd_sc_hd__a21oi_1 _10667_ (.A1(_04127_),
    .A2(_04795_),
    .B1(net3726),
    .Y(_04798_));
 sky130_fd_sc_hd__a31o_1 _10668_ (.A1(net3726),
    .A2(_04127_),
    .A3(_04795_),
    .B1(_00228_),
    .X(_04799_));
 sky130_fd_sc_hd__nor2_1 _10669_ (.A(_04798_),
    .B(_04799_),
    .Y(_00161_));
 sky130_fd_sc_hd__and3_1 _10670_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .B(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .C(_04373_),
    .X(_04800_));
 sky130_fd_sc_hd__a31o_1 _10671_ (.A1(net3330),
    .A2(_04355_),
    .A3(_04800_),
    .B1(\c.genblk1.genblk1.subs.c0.cfgd ),
    .X(_04801_));
 sky130_fd_sc_hd__and2_1 _10672_ (.A(_00196_),
    .B(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__clkbuf_1 _10673_ (.A(_04802_),
    .X(_00162_));
 sky130_fd_sc_hd__and3b_1 _10674_ (.A_N(_04800_),
    .B(_04355_),
    .C(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(_04803_));
 sky130_fd_sc_hd__nor2_1 _10675_ (.A(_00268_),
    .B(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__o21a_1 _10676_ (.A1(net3270),
    .A2(_04355_),
    .B1(_04804_),
    .X(_00163_));
 sky130_fd_sc_hd__and2_1 _10677_ (.A(net3275),
    .B(_04803_),
    .X(_04805_));
 sky130_fd_sc_hd__a21oi_1 _10678_ (.A1(net3270),
    .A2(_04355_),
    .B1(net3275),
    .Y(_04806_));
 sky130_fd_sc_hd__nor3_1 _10679_ (.A(_04531_),
    .B(_04805_),
    .C(_04806_),
    .Y(_00164_));
 sky130_fd_sc_hd__and3_1 _10680_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .B(net3275),
    .C(_04803_),
    .X(_04807_));
 sky130_fd_sc_hd__nor2_1 _10681_ (.A(_00268_),
    .B(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hd__o21a_1 _10682_ (.A1(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .A2(_04805_),
    .B1(_04808_),
    .X(_00165_));
 sky130_fd_sc_hd__a21oi_1 _10683_ (.A1(_04345_),
    .A2(_04807_),
    .B1(_04729_),
    .Y(_04809_));
 sky130_fd_sc_hd__o21a_1 _10684_ (.A1(_04345_),
    .A2(_04807_),
    .B1(_04809_),
    .X(_00166_));
 sky130_fd_sc_hd__a21oi_1 _10685_ (.A1(_04345_),
    .A2(_04807_),
    .B1(net3831),
    .Y(_04810_));
 sky130_fd_sc_hd__and3_1 _10686_ (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .B(_04345_),
    .C(_04807_),
    .X(_04811_));
 sky130_fd_sc_hd__nor3_1 _10687_ (.A(_04531_),
    .B(_04810_),
    .C(_04811_),
    .Y(_00167_));
 sky130_fd_sc_hd__a21oi_1 _10688_ (.A1(net3728),
    .A2(_04811_),
    .B1(_04520_),
    .Y(_04812_));
 sky130_fd_sc_hd__o21a_1 _10689_ (.A1(net3728),
    .A2(_04811_),
    .B1(_04812_),
    .X(_00168_));
 sky130_fd_sc_hd__or3_1 _10690_ (.A(_02759_),
    .B(_00793_),
    .C(_03993_),
    .X(_04813_));
 sky130_fd_sc_hd__o21a_1 _10691_ (.A1(net3846),
    .A2(_02525_),
    .B1(_04813_),
    .X(_00169_));
 sky130_fd_sc_hd__dfxtp_1 _10692_ (.CLK(clknet_leaf_29_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10693_ (.CLK(clknet_leaf_28_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10694_ (.CLK(clknet_leaf_30_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10695_ (.CLK(clknet_leaf_29_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10696_ (.CLK(clknet_leaf_71_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10697_ (.CLK(clknet_leaf_72_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10698_ (.CLK(clknet_leaf_71_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10699_ (.CLK(clknet_leaf_68_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10700_ (.CLK(clknet_leaf_65_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10701_ (.CLK(clknet_leaf_71_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10702_ (.CLK(clknet_leaf_73_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10703_ (.CLK(clknet_leaf_71_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10704_ (.CLK(clknet_leaf_65_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10705_ (.CLK(clknet_leaf_72_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10706_ (.CLK(clknet_leaf_65_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10707_ (.CLK(clknet_leaf_71_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10708_ (.CLK(clknet_leaf_66_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10709_ (.CLK(clknet_leaf_67_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10710_ (.CLK(clknet_leaf_66_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10711_ (.CLK(clknet_leaf_66_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10712_ (.CLK(clknet_leaf_71_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10713_ (.CLK(clknet_leaf_72_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10714_ (.CLK(clknet_leaf_73_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10715_ (.CLK(clknet_leaf_66_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10716_ (.CLK(clknet_leaf_73_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10717_ (.CLK(clknet_leaf_72_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10718_ (.CLK(clknet_leaf_72_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10719_ (.CLK(clknet_leaf_68_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10720_ (.CLK(clknet_leaf_73_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10721_ (.CLK(clknet_leaf_72_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10722_ (.CLK(clknet_leaf_73_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _10723_ (.CLK(clknet_leaf_66_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _10724_ (.CLK(clknet_leaf_64_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _10725_ (.CLK(clknet_leaf_65_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _10726_ (.CLK(clknet_leaf_64_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _10727_ (.CLK(clknet_leaf_64_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _10728_ (.CLK(clknet_leaf_65_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _10729_ (.CLK(clknet_leaf_31_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _10730_ (.CLK(clknet_leaf_29_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _10731_ (.CLK(clknet_leaf_29_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _10732_ (.CLK(clknet_leaf_28_clk),
    .D(net497),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10733_ (.CLK(clknet_leaf_28_clk),
    .D(net1556),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10734_ (.CLK(clknet_leaf_29_clk),
    .D(net605),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10735_ (.CLK(clknet_leaf_29_clk),
    .D(net2372),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10736_ (.CLK(clknet_leaf_71_clk),
    .D(net1283),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10737_ (.CLK(clknet_leaf_71_clk),
    .D(net588),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10738_ (.CLK(clknet_leaf_71_clk),
    .D(net1136),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10739_ (.CLK(clknet_leaf_68_clk),
    .D(net2860),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10740_ (.CLK(clknet_leaf_65_clk),
    .D(net2276),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10741_ (.CLK(clknet_leaf_74_clk),
    .D(net414),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10742_ (.CLK(clknet_leaf_73_clk),
    .D(net2342),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10743_ (.CLK(clknet_leaf_71_clk),
    .D(net1514),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10744_ (.CLK(clknet_leaf_65_clk),
    .D(net2212),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10745_ (.CLK(clknet_leaf_72_clk),
    .D(net2602),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10746_ (.CLK(clknet_leaf_65_clk),
    .D(net2328),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10747_ (.CLK(clknet_leaf_70_clk),
    .D(net423),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10748_ (.CLK(clknet_leaf_66_clk),
    .D(net877),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10749_ (.CLK(clknet_leaf_67_clk),
    .D(net2566),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10750_ (.CLK(clknet_leaf_66_clk),
    .D(net1065),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10751_ (.CLK(clknet_leaf_66_clk),
    .D(net892),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10752_ (.CLK(clknet_leaf_71_clk),
    .D(net2104),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10753_ (.CLK(clknet_leaf_73_clk),
    .D(net359),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10754_ (.CLK(clknet_leaf_73_clk),
    .D(net2415),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10755_ (.CLK(clknet_leaf_66_clk),
    .D(net838),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10756_ (.CLK(clknet_leaf_73_clk),
    .D(net1669),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10757_ (.CLK(clknet_leaf_72_clk),
    .D(net2246),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10758_ (.CLK(clknet_leaf_73_clk),
    .D(net442),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10759_ (.CLK(clknet_leaf_70_clk),
    .D(net56),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10760_ (.CLK(clknet_leaf_73_clk),
    .D(net2801),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10761_ (.CLK(clknet_leaf_73_clk),
    .D(net666),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10762_ (.CLK(clknet_leaf_73_clk),
    .D(net2838),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _10763_ (.CLK(clknet_leaf_71_clk),
    .D(net46),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _10764_ (.CLK(clknet_leaf_64_clk),
    .D(net1756),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _10765_ (.CLK(clknet_leaf_65_clk),
    .D(net1715),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _10766_ (.CLK(clknet_leaf_63_clk),
    .D(net425),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _10767_ (.CLK(clknet_leaf_64_clk),
    .D(net1036),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _10768_ (.CLK(clknet_leaf_65_clk),
    .D(net2495),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _10769_ (.CLK(clknet_leaf_29_clk),
    .D(net260),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _10770_ (.CLK(clknet_leaf_29_clk),
    .D(net1457),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _10771_ (.CLK(clknet_leaf_29_clk),
    .D(net1837),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _10772_ (.CLK(clknet_leaf_28_clk),
    .D(net2701),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10773_ (.CLK(clknet_leaf_28_clk),
    .D(net2671),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10774_ (.CLK(clknet_leaf_30_clk),
    .D(net487),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10775_ (.CLK(clknet_leaf_29_clk),
    .D(net2046),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10776_ (.CLK(clknet_leaf_71_clk),
    .D(net1577),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10777_ (.CLK(clknet_leaf_71_clk),
    .D(net1639),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10778_ (.CLK(clknet_leaf_71_clk),
    .D(net1506),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10779_ (.CLK(clknet_leaf_68_clk),
    .D(net2642),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10780_ (.CLK(clknet_leaf_65_clk),
    .D(net2345),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10781_ (.CLK(clknet_leaf_74_clk),
    .D(net2028),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10782_ (.CLK(clknet_leaf_74_clk),
    .D(net756),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10783_ (.CLK(clknet_leaf_71_clk),
    .D(net2649),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10784_ (.CLK(clknet_leaf_67_clk),
    .D(net332),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10785_ (.CLK(clknet_leaf_72_clk),
    .D(net1684),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10786_ (.CLK(clknet_leaf_65_clk),
    .D(net1867),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10787_ (.CLK(clknet_leaf_70_clk),
    .D(net1390),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10788_ (.CLK(clknet_leaf_72_clk),
    .D(net49),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10789_ (.CLK(clknet_leaf_67_clk),
    .D(net2161),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10790_ (.CLK(clknet_leaf_66_clk),
    .D(net841),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10791_ (.CLK(clknet_leaf_72_clk),
    .D(net47),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10792_ (.CLK(clknet_leaf_73_clk),
    .D(net389),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10793_ (.CLK(clknet_leaf_73_clk),
    .D(net1970),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10794_ (.CLK(clknet_leaf_73_clk),
    .D(net2472),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10795_ (.CLK(clknet_leaf_72_clk),
    .D(net48),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10796_ (.CLK(clknet_leaf_73_clk),
    .D(net1356),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10797_ (.CLK(clknet_leaf_72_clk),
    .D(net2901),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10798_ (.CLK(clknet_leaf_73_clk),
    .D(net1908),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10799_ (.CLK(clknet_leaf_70_clk),
    .D(net1386),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10800_ (.CLK(clknet_leaf_73_clk),
    .D(net2807),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10801_ (.CLK(clknet_leaf_72_clk),
    .D(net622),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10802_ (.CLK(clknet_leaf_73_clk),
    .D(net2863),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _10803_ (.CLK(clknet_leaf_71_clk),
    .D(net2087),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _10804_ (.CLK(clknet_leaf_63_clk),
    .D(net443),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _10805_ (.CLK(clknet_leaf_67_clk),
    .D(net495),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _10806_ (.CLK(clknet_leaf_65_clk),
    .D(net158),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _10807_ (.CLK(clknet_leaf_64_clk),
    .D(net1819),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _10808_ (.CLK(clknet_leaf_65_clk),
    .D(net1903),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _10809_ (.CLK(clknet_leaf_29_clk),
    .D(net1501),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _10810_ (.CLK(clknet_leaf_65_clk),
    .D(net520),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _10811_ (.CLK(clknet_leaf_65_clk),
    .D(net550),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_2 _10812_ (.CLK(clknet_leaf_28_clk),
    .D(net1023),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[0] ));
 sky130_fd_sc_hd__dfxtp_2 _10813_ (.CLK(clknet_leaf_65_clk),
    .D(net593),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10814_ (.CLK(clknet_leaf_64_clk),
    .D(net293),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _10815_ (.CLK(clknet_leaf_29_clk),
    .D(net1154),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[3] ));
 sky130_fd_sc_hd__dfxtp_2 _10816_ (.CLK(clknet_leaf_71_clk),
    .D(net1519),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[4] ));
 sky130_fd_sc_hd__dfxtp_4 _10817_ (.CLK(clknet_leaf_71_clk),
    .D(net1048),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ));
 sky130_fd_sc_hd__dfxtp_2 _10818_ (.CLK(clknet_leaf_74_clk),
    .D(net441),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _10819_ (.CLK(clknet_leaf_69_clk),
    .D(net58),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _10820_ (.CLK(clknet_leaf_65_clk),
    .D(net1702),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _10821_ (.CLK(clknet_leaf_74_clk),
    .D(net2596),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[9] ));
 sky130_fd_sc_hd__dfxtp_4 _10822_ (.CLK(clknet_leaf_74_clk),
    .D(net1078),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ));
 sky130_fd_sc_hd__dfxtp_2 _10823_ (.CLK(clknet_leaf_71_clk),
    .D(net1536),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _10824_ (.CLK(clknet_leaf_67_clk),
    .D(net1412),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _10825_ (.CLK(clknet_leaf_72_clk),
    .D(net2484),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _10826_ (.CLK(clknet_leaf_67_clk),
    .D(net335),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[14] ));
 sky130_fd_sc_hd__dfxtp_4 _10827_ (.CLK(clknet_leaf_71_clk),
    .D(net482),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _10828_ (.CLK(clknet_leaf_71_clk),
    .D(net384),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[16] ));
 sky130_fd_sc_hd__dfxtp_1 _10829_ (.CLK(clknet_leaf_66_clk),
    .D(net943),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[17] ));
 sky130_fd_sc_hd__dfxtp_1 _10830_ (.CLK(clknet_leaf_66_clk),
    .D(net1781),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[18] ));
 sky130_fd_sc_hd__dfxtp_1 _10831_ (.CLK(clknet_leaf_72_clk),
    .D(net1966),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[19] ));
 sky130_fd_sc_hd__dfxtp_4 _10832_ (.CLK(clknet_leaf_74_clk),
    .D(net413),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ));
 sky130_fd_sc_hd__dfxtp_2 _10833_ (.CLK(clknet_leaf_73_clk),
    .D(net2253),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ));
 sky130_fd_sc_hd__dfxtp_1 _10834_ (.CLK(clknet_leaf_73_clk),
    .D(net2604),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _10835_ (.CLK(clknet_leaf_72_clk),
    .D(net1842),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[23] ));
 sky130_fd_sc_hd__dfxtp_1 _10836_ (.CLK(clknet_leaf_75_clk),
    .D(net746),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[24] ));
 sky130_fd_sc_hd__dfxtp_2 _10837_ (.CLK(clknet_leaf_72_clk),
    .D(net1604),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ));
 sky130_fd_sc_hd__dfxtp_2 _10838_ (.CLK(clknet_leaf_73_clk),
    .D(net2007),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ));
 sky130_fd_sc_hd__dfxtp_1 _10839_ (.CLK(clknet_leaf_70_clk),
    .D(net2309),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[27] ));
 sky130_fd_sc_hd__dfxtp_1 _10840_ (.CLK(clknet_leaf_75_clk),
    .D(net731),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[28] ));
 sky130_fd_sc_hd__dfxtp_1 _10841_ (.CLK(clknet_leaf_72_clk),
    .D(net1933),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[29] ));
 sky130_fd_sc_hd__dfxtp_4 _10842_ (.CLK(clknet_leaf_75_clk),
    .D(net714),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ));
 sky130_fd_sc_hd__dfxtp_2 _10843_ (.CLK(clknet_leaf_72_clk),
    .D(net437),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ));
 sky130_fd_sc_hd__dfxtp_1 _10844_ (.CLK(clknet_leaf_63_clk),
    .D(net1589),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[32] ));
 sky130_fd_sc_hd__dfxtp_1 _10845_ (.CLK(clknet_leaf_67_clk),
    .D(net1948),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[33] ));
 sky130_fd_sc_hd__dfxtp_1 _10846_ (.CLK(clknet_leaf_63_clk),
    .D(net266),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[34] ));
 sky130_fd_sc_hd__dfxtp_2 _10847_ (.CLK(clknet_leaf_64_clk),
    .D(net1024),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[35] ));
 sky130_fd_sc_hd__dfxtp_2 _10848_ (.CLK(clknet_leaf_65_clk),
    .D(net983),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[36] ));
 sky130_fd_sc_hd__dfxtp_1 _10849_ (.CLK(clknet_leaf_30_clk),
    .D(net543),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[37] ));
 sky130_fd_sc_hd__dfxtp_1 _10850_ (.CLK(clknet_leaf_65_clk),
    .D(net2610),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[38] ));
 sky130_fd_sc_hd__dfxtp_1 _10851_ (.CLK(clknet_leaf_65_clk),
    .D(net1554),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[39] ));
 sky130_fd_sc_hd__dfxtp_1 _10852_ (.CLK(clknet_leaf_67_clk),
    .D(_00016_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _10853_ (.CLK(clknet_leaf_68_clk),
    .D(_00017_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _10854_ (.CLK(clknet_leaf_68_clk),
    .D(_00018_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10855_ (.CLK(clknet_leaf_68_clk),
    .D(_00019_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _10856_ (.CLK(clknet_leaf_67_clk),
    .D(_00020_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _10857_ (.CLK(clknet_leaf_66_clk),
    .D(_00021_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _10858_ (.CLK(clknet_leaf_67_clk),
    .D(_00022_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _10859_ (.CLK(clknet_leaf_64_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__dfxtp_2 _10860_ (.CLK(clknet_leaf_43_clk),
    .D(net3620),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__dfxtp_2 _10861_ (.CLK(clknet_leaf_55_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__dfxtp_2 _10862_ (.CLK(clknet_leaf_30_clk),
    .D(net3679),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__dfxtp_4 _10863_ (.CLK(clknet_leaf_43_clk),
    .D(net3702),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__dfxtp_4 _10864_ (.CLK(clknet_leaf_43_clk),
    .D(net3577),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__dfxtp_4 _10865_ (.CLK(clknet_leaf_64_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__dfxtp_4 _10866_ (.CLK(clknet_leaf_42_clk),
    .D(net3844),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _10867_ (.CLK(clknet_leaf_29_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10868_ (.CLK(clknet_leaf_29_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10869_ (.CLK(clknet_leaf_30_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10870_ (.CLK(clknet_leaf_30_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10871_ (.CLK(clknet_leaf_40_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10872_ (.CLK(clknet_leaf_45_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10873_ (.CLK(clknet_leaf_45_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10874_ (.CLK(clknet_leaf_45_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10875_ (.CLK(clknet_leaf_45_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10876_ (.CLK(clknet_leaf_46_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10877_ (.CLK(clknet_leaf_45_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10878_ (.CLK(clknet_leaf_45_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10879_ (.CLK(clknet_leaf_43_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10880_ (.CLK(clknet_leaf_43_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10881_ (.CLK(clknet_leaf_43_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10882_ (.CLK(clknet_leaf_43_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10883_ (.CLK(clknet_leaf_42_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10884_ (.CLK(clknet_leaf_41_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10885_ (.CLK(clknet_leaf_42_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10886_ (.CLK(clknet_leaf_42_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10887_ (.CLK(clknet_leaf_44_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10888_ (.CLK(clknet_leaf_46_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10889_ (.CLK(clknet_leaf_44_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10890_ (.CLK(clknet_leaf_46_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10891_ (.CLK(clknet_leaf_46_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10892_ (.CLK(clknet_leaf_47_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10893_ (.CLK(clknet_leaf_46_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10894_ (.CLK(clknet_leaf_46_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10895_ (.CLK(clknet_leaf_47_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10896_ (.CLK(clknet_leaf_46_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10897_ (.CLK(clknet_leaf_44_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _10898_ (.CLK(clknet_leaf_45_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _10899_ (.CLK(clknet_leaf_30_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _10900_ (.CLK(clknet_leaf_30_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _10901_ (.CLK(clknet_leaf_30_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _10902_ (.CLK(clknet_leaf_42_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _10903_ (.CLK(clknet_leaf_40_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _10904_ (.CLK(clknet_leaf_39_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _10905_ (.CLK(clknet_leaf_40_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _10906_ (.CLK(clknet_leaf_39_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _10907_ (.CLK(clknet_leaf_31_clk),
    .D(net109),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10908_ (.CLK(clknet_leaf_30_clk),
    .D(net558),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10909_ (.CLK(clknet_leaf_30_clk),
    .D(net1598),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10910_ (.CLK(clknet_leaf_30_clk),
    .D(net2094),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10911_ (.CLK(clknet_leaf_40_clk),
    .D(net1435),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10912_ (.CLK(clknet_leaf_45_clk),
    .D(net1761),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10913_ (.CLK(clknet_leaf_45_clk),
    .D(net2401),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10914_ (.CLK(clknet_leaf_45_clk),
    .D(net2379),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10915_ (.CLK(clknet_leaf_45_clk),
    .D(net1662),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10916_ (.CLK(clknet_leaf_46_clk),
    .D(net2355),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10917_ (.CLK(clknet_leaf_46_clk),
    .D(net689),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10918_ (.CLK(clknet_leaf_45_clk),
    .D(net2751),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10919_ (.CLK(clknet_leaf_43_clk),
    .D(net2251),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10920_ (.CLK(clknet_leaf_43_clk),
    .D(net2612),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10921_ (.CLK(clknet_leaf_43_clk),
    .D(net2392),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10922_ (.CLK(clknet_leaf_43_clk),
    .D(net1606),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10923_ (.CLK(clknet_leaf_42_clk),
    .D(net1218),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10924_ (.CLK(clknet_leaf_41_clk),
    .D(net2655),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10925_ (.CLK(clknet_leaf_42_clk),
    .D(net1782),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10926_ (.CLK(clknet_leaf_42_clk),
    .D(net1442),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10927_ (.CLK(clknet_leaf_44_clk),
    .D(net1015),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10928_ (.CLK(clknet_leaf_46_clk),
    .D(net2710),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10929_ (.CLK(clknet_leaf_44_clk),
    .D(net1063),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10930_ (.CLK(clknet_leaf_46_clk),
    .D(net2845),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10931_ (.CLK(clknet_leaf_46_clk),
    .D(net2231),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10932_ (.CLK(clknet_leaf_47_clk),
    .D(net2006),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10933_ (.CLK(clknet_leaf_46_clk),
    .D(net2219),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10934_ (.CLK(clknet_leaf_47_clk),
    .D(net313),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10935_ (.CLK(clknet_leaf_47_clk),
    .D(net2707),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10936_ (.CLK(clknet_leaf_46_clk),
    .D(net2916),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10937_ (.CLK(clknet_leaf_44_clk),
    .D(net1072),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _10938_ (.CLK(clknet_leaf_46_clk),
    .D(net708),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _10939_ (.CLK(clknet_leaf_30_clk),
    .D(net2519),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _10940_ (.CLK(clknet_leaf_30_clk),
    .D(net2629),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _10941_ (.CLK(clknet_leaf_30_clk),
    .D(net2639),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _10942_ (.CLK(clknet_leaf_31_clk),
    .D(net296),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _10943_ (.CLK(clknet_leaf_40_clk),
    .D(net1391),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _10944_ (.CLK(clknet_leaf_39_clk),
    .D(net1635),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _10945_ (.CLK(clknet_leaf_40_clk),
    .D(net1573),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _10946_ (.CLK(clknet_leaf_40_clk),
    .D(net797),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _10947_ (.CLK(clknet_leaf_31_clk),
    .D(net1287),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10948_ (.CLK(clknet_leaf_29_clk),
    .D(net650),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10949_ (.CLK(clknet_leaf_30_clk),
    .D(net2209),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10950_ (.CLK(clknet_leaf_30_clk),
    .D(net2195),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10951_ (.CLK(clknet_leaf_40_clk),
    .D(net2183),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10952_ (.CLK(clknet_leaf_45_clk),
    .D(net2508),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10953_ (.CLK(clknet_leaf_45_clk),
    .D(net1717),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10954_ (.CLK(clknet_leaf_45_clk),
    .D(net1521),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10955_ (.CLK(clknet_leaf_45_clk),
    .D(net1086),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10956_ (.CLK(clknet_leaf_46_clk),
    .D(net2623),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10957_ (.CLK(clknet_leaf_46_clk),
    .D(net1082),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10958_ (.CLK(clknet_leaf_45_clk),
    .D(net1783),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10959_ (.CLK(clknet_leaf_43_clk),
    .D(net907),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10960_ (.CLK(clknet_leaf_43_clk),
    .D(net1912),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10961_ (.CLK(clknet_leaf_43_clk),
    .D(net910),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10962_ (.CLK(clknet_leaf_43_clk),
    .D(net1998),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10963_ (.CLK(clknet_leaf_42_clk),
    .D(net1004),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10964_ (.CLK(clknet_leaf_41_clk),
    .D(net1929),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10965_ (.CLK(clknet_leaf_42_clk),
    .D(net1387),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10966_ (.CLK(clknet_leaf_42_clk),
    .D(net2045),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10967_ (.CLK(clknet_leaf_44_clk),
    .D(net872),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10968_ (.CLK(clknet_leaf_46_clk),
    .D(net1984),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10969_ (.CLK(clknet_leaf_44_clk),
    .D(net966),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10970_ (.CLK(clknet_leaf_46_clk),
    .D(net2126),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10971_ (.CLK(clknet_leaf_46_clk),
    .D(net2337),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10972_ (.CLK(clknet_leaf_47_clk),
    .D(net1887),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10973_ (.CLK(clknet_leaf_46_clk),
    .D(net2116),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10974_ (.CLK(clknet_leaf_47_clk),
    .D(net1713),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10975_ (.CLK(clknet_leaf_47_clk),
    .D(net1541),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10976_ (.CLK(clknet_leaf_47_clk),
    .D(net331),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10977_ (.CLK(clknet_leaf_43_clk),
    .D(net312),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _10978_ (.CLK(clknet_leaf_45_clk),
    .D(net481),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _10979_ (.CLK(clknet_leaf_31_clk),
    .D(net107),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _10980_ (.CLK(clknet_leaf_30_clk),
    .D(net2021),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _10981_ (.CLK(clknet_leaf_30_clk),
    .D(net2723),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _10982_ (.CLK(clknet_leaf_42_clk),
    .D(net769),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _10983_ (.CLK(clknet_leaf_40_clk),
    .D(net992),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _10984_ (.CLK(clknet_leaf_39_clk),
    .D(net1246),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _10985_ (.CLK(clknet_leaf_45_clk),
    .D(net174),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _10986_ (.CLK(clknet_leaf_40_clk),
    .D(net885),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_2 _10987_ (.CLK(clknet_leaf_29_clk),
    .D(net230),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[0] ));
 sky130_fd_sc_hd__dfxtp_2 _10988_ (.CLK(clknet_leaf_30_clk),
    .D(net455),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10989_ (.CLK(clknet_leaf_64_clk),
    .D(net317),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _10990_ (.CLK(clknet_leaf_30_clk),
    .D(net1829),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _10991_ (.CLK(clknet_leaf_40_clk),
    .D(net1210),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[4] ));
 sky130_fd_sc_hd__dfxtp_4 _10992_ (.CLK(clknet_leaf_45_clk),
    .D(net1123),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ));
 sky130_fd_sc_hd__dfxtp_4 _10993_ (.CLK(clknet_leaf_45_clk),
    .D(net866),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _10994_ (.CLK(clknet_leaf_45_clk),
    .D(net1613),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _10995_ (.CLK(clknet_leaf_44_clk),
    .D(net803),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _10996_ (.CLK(clknet_leaf_46_clk),
    .D(net2815),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[9] ));
 sky130_fd_sc_hd__dfxtp_4 _10997_ (.CLK(clknet_leaf_45_clk),
    .D(net349),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ));
 sky130_fd_sc_hd__dfxtp_4 _10998_ (.CLK(clknet_leaf_45_clk),
    .D(net1300),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _10999_ (.CLK(clknet_leaf_43_clk),
    .D(net1186),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _11000_ (.CLK(clknet_leaf_55_clk),
    .D(net510),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _11001_ (.CLK(clknet_leaf_55_clk),
    .D(net294),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[14] ));
 sky130_fd_sc_hd__dfxtp_2 _11002_ (.CLK(clknet_leaf_43_clk),
    .D(net1032),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _11003_ (.CLK(clknet_leaf_42_clk),
    .D(net921),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ));
 sky130_fd_sc_hd__dfxtp_1 _11004_ (.CLK(clknet_leaf_42_clk),
    .D(net738),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[17] ));
 sky130_fd_sc_hd__dfxtp_1 _11005_ (.CLK(clknet_leaf_42_clk),
    .D(net1576),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[18] ));
 sky130_fd_sc_hd__dfxtp_1 _11006_ (.CLK(clknet_leaf_42_clk),
    .D(net1235),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[19] ));
 sky130_fd_sc_hd__dfxtp_2 _11007_ (.CLK(clknet_leaf_44_clk),
    .D(net865),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[20] ));
 sky130_fd_sc_hd__dfxtp_2 _11008_ (.CLK(clknet_leaf_46_clk),
    .D(net998),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ));
 sky130_fd_sc_hd__dfxtp_1 _11009_ (.CLK(clknet_leaf_44_clk),
    .D(net906),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _11010_ (.CLK(clknet_leaf_46_clk),
    .D(net1934),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[23] ));
 sky130_fd_sc_hd__dfxtp_1 _11011_ (.CLK(clknet_leaf_46_clk),
    .D(net2853),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[24] ));
 sky130_fd_sc_hd__dfxtp_2 _11012_ (.CLK(clknet_leaf_47_clk),
    .D(net1384),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[25] ));
 sky130_fd_sc_hd__dfxtp_2 _11013_ (.CLK(clknet_leaf_47_clk),
    .D(net315),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ));
 sky130_fd_sc_hd__dfxtp_1 _11014_ (.CLK(clknet_leaf_47_clk),
    .D(net1396),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[27] ));
 sky130_fd_sc_hd__dfxtp_1 _11015_ (.CLK(clknet_leaf_47_clk),
    .D(net2854),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[28] ));
 sky130_fd_sc_hd__dfxtp_1 _11016_ (.CLK(clknet_leaf_47_clk),
    .D(net1802),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[29] ));
 sky130_fd_sc_hd__dfxtp_2 _11017_ (.CLK(clknet_leaf_43_clk),
    .D(net2929),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[30] ));
 sky130_fd_sc_hd__dfxtp_2 _11018_ (.CLK(clknet_leaf_44_clk),
    .D(net807),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ));
 sky130_fd_sc_hd__dfxtp_1 _11019_ (.CLK(clknet_leaf_31_clk),
    .D(net1923),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[32] ));
 sky130_fd_sc_hd__dfxtp_1 _11020_ (.CLK(clknet_leaf_30_clk),
    .D(net1335),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[33] ));
 sky130_fd_sc_hd__dfxtp_1 _11021_ (.CLK(clknet_leaf_30_clk),
    .D(net2855),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[34] ));
 sky130_fd_sc_hd__dfxtp_2 _11022_ (.CLK(clknet_leaf_30_clk),
    .D(net196),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[35] ));
 sky130_fd_sc_hd__dfxtp_2 _11023_ (.CLK(clknet_leaf_40_clk),
    .D(net923),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ));
 sky130_fd_sc_hd__dfxtp_2 _11024_ (.CLK(clknet_leaf_40_clk),
    .D(net773),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[37] ));
 sky130_fd_sc_hd__dfxtp_1 _11025_ (.CLK(clknet_leaf_45_clk),
    .D(net1660),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ));
 sky130_fd_sc_hd__dfxtp_1 _11026_ (.CLK(clknet_leaf_40_clk),
    .D(net1777),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[39] ));
 sky130_fd_sc_hd__dfxtp_1 _11027_ (.CLK(clknet_leaf_42_clk),
    .D(_00023_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _11028_ (.CLK(clknet_leaf_42_clk),
    .D(_00024_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11029_ (.CLK(clknet_leaf_42_clk),
    .D(_00025_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11030_ (.CLK(clknet_leaf_43_clk),
    .D(_00026_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11031_ (.CLK(clknet_leaf_44_clk),
    .D(_00027_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11032_ (.CLK(clknet_leaf_44_clk),
    .D(_00028_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11033_ (.CLK(clknet_leaf_41_clk),
    .D(_00029_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _11034_ (.CLK(clknet_leaf_63_clk),
    .D(net3745),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__dfxtp_4 _11035_ (.CLK(clknet_leaf_55_clk),
    .D(net3424),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__dfxtp_4 _11036_ (.CLK(clknet_leaf_53_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__dfxtp_4 _11037_ (.CLK(clknet_leaf_63_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__dfxtp_4 _11038_ (.CLK(clknet_leaf_56_clk),
    .D(net4226),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__dfxtp_4 _11039_ (.CLK(clknet_leaf_59_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__dfxtp_4 _11040_ (.CLK(clknet_leaf_56_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__dfxtp_4 _11041_ (.CLK(clknet_leaf_55_clk),
    .D(net3506),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11042_ (.CLK(clknet_leaf_64_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11043_ (.CLK(clknet_leaf_64_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11044_ (.CLK(clknet_leaf_64_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11045_ (.CLK(clknet_leaf_63_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11046_ (.CLK(clknet_leaf_55_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11047_ (.CLK(clknet_leaf_48_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11048_ (.CLK(clknet_leaf_47_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11049_ (.CLK(clknet_leaf_47_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11050_ (.CLK(clknet_leaf_44_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11051_ (.CLK(clknet_leaf_48_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11052_ (.CLK(clknet_leaf_48_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11053_ (.CLK(clknet_leaf_50_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11054_ (.CLK(clknet_leaf_51_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11055_ (.CLK(clknet_leaf_51_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11056_ (.CLK(clknet_leaf_52_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11057_ (.CLK(clknet_leaf_56_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11058_ (.CLK(clknet_leaf_56_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11059_ (.CLK(clknet_leaf_56_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11060_ (.CLK(clknet_leaf_56_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11061_ (.CLK(clknet_leaf_56_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11062_ (.CLK(clknet_leaf_58_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11063_ (.CLK(clknet_leaf_57_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11064_ (.CLK(clknet_leaf_57_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11065_ (.CLK(clknet_leaf_57_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11066_ (.CLK(clknet_leaf_58_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11067_ (.CLK(clknet_leaf_59_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11068_ (.CLK(clknet_leaf_57_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11069_ (.CLK(clknet_leaf_59_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11070_ (.CLK(clknet_leaf_59_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11071_ (.CLK(clknet_leaf_59_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11072_ (.CLK(clknet_leaf_53_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11073_ (.CLK(clknet_leaf_52_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11074_ (.CLK(clknet_leaf_48_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11075_ (.CLK(clknet_leaf_48_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11076_ (.CLK(clknet_leaf_48_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11077_ (.CLK(clknet_leaf_48_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11078_ (.CLK(clknet_leaf_55_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11079_ (.CLK(clknet_leaf_53_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11080_ (.CLK(clknet_leaf_54_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11081_ (.CLK(clknet_leaf_53_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _11082_ (.CLK(clknet_leaf_64_clk),
    .D(net1680),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11083_ (.CLK(clknet_leaf_55_clk),
    .D(net794),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11084_ (.CLK(clknet_leaf_64_clk),
    .D(net1626),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11085_ (.CLK(clknet_leaf_63_clk),
    .D(net1370),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11086_ (.CLK(clknet_leaf_55_clk),
    .D(net1409),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11087_ (.CLK(clknet_leaf_48_clk),
    .D(net2740),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11088_ (.CLK(clknet_leaf_47_clk),
    .D(net2010),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11089_ (.CLK(clknet_leaf_47_clk),
    .D(net1339),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11090_ (.CLK(clknet_leaf_54_clk),
    .D(net817),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11091_ (.CLK(clknet_leaf_48_clk),
    .D(net2788),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11092_ (.CLK(clknet_leaf_48_clk),
    .D(net1336),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11093_ (.CLK(clknet_leaf_50_clk),
    .D(net2453),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11094_ (.CLK(clknet_leaf_51_clk),
    .D(net2605),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11095_ (.CLK(clknet_leaf_51_clk),
    .D(net2143),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11096_ (.CLK(clknet_leaf_52_clk),
    .D(net1363),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11097_ (.CLK(clknet_leaf_56_clk),
    .D(net1567),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11098_ (.CLK(clknet_leaf_56_clk),
    .D(net1564),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11099_ (.CLK(clknet_leaf_56_clk),
    .D(net1066),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11100_ (.CLK(clknet_leaf_56_clk),
    .D(net2675),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11101_ (.CLK(clknet_leaf_63_clk),
    .D(net363),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11102_ (.CLK(clknet_leaf_58_clk),
    .D(net1144),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11103_ (.CLK(clknet_leaf_57_clk),
    .D(net1088),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11104_ (.CLK(clknet_leaf_57_clk),
    .D(net1085),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11105_ (.CLK(clknet_leaf_56_clk),
    .D(net356),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11106_ (.CLK(clknet_leaf_58_clk),
    .D(net2142),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11107_ (.CLK(clknet_leaf_59_clk),
    .D(net1448),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11108_ (.CLK(clknet_leaf_57_clk),
    .D(net913),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11109_ (.CLK(clknet_leaf_59_clk),
    .D(net1655),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11110_ (.CLK(clknet_leaf_59_clk),
    .D(net2530),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11111_ (.CLK(clknet_leaf_59_clk),
    .D(net1875),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11112_ (.CLK(clknet_leaf_53_clk),
    .D(net890),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11113_ (.CLK(clknet_leaf_52_clk),
    .D(net928),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11114_ (.CLK(clknet_leaf_48_clk),
    .D(net2174),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11115_ (.CLK(clknet_leaf_48_clk),
    .D(net1938),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11116_ (.CLK(clknet_leaf_48_clk),
    .D(net2480),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11117_ (.CLK(clknet_leaf_48_clk),
    .D(net2466),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11118_ (.CLK(clknet_leaf_54_clk),
    .D(net128),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11119_ (.CLK(clknet_leaf_53_clk),
    .D(net816),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11120_ (.CLK(clknet_leaf_54_clk),
    .D(net811),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11121_ (.CLK(clknet_leaf_54_clk),
    .D(net696),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _11122_ (.CLK(clknet_leaf_64_clk),
    .D(net2650),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11123_ (.CLK(clknet_leaf_55_clk),
    .D(net843),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11124_ (.CLK(clknet_leaf_64_clk),
    .D(net2780),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11125_ (.CLK(clknet_leaf_63_clk),
    .D(net1892),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11126_ (.CLK(clknet_leaf_55_clk),
    .D(net1141),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11127_ (.CLK(clknet_leaf_47_clk),
    .D(net718),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11128_ (.CLK(clknet_leaf_47_clk),
    .D(net2118),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11129_ (.CLK(clknet_leaf_44_clk),
    .D(net914),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11130_ (.CLK(clknet_leaf_54_clk),
    .D(net820),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11131_ (.CLK(clknet_leaf_47_clk),
    .D(net614),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11132_ (.CLK(clknet_leaf_48_clk),
    .D(net2783),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11133_ (.CLK(clknet_leaf_50_clk),
    .D(net1883),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11134_ (.CLK(clknet_leaf_51_clk),
    .D(net1663),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11135_ (.CLK(clknet_leaf_51_clk),
    .D(net1096),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11136_ (.CLK(clknet_leaf_52_clk),
    .D(net1101),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11137_ (.CLK(clknet_leaf_56_clk),
    .D(net2488),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11138_ (.CLK(clknet_leaf_56_clk),
    .D(net2479),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11139_ (.CLK(clknet_leaf_63_clk),
    .D(net383),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11140_ (.CLK(clknet_leaf_56_clk),
    .D(net1142),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11141_ (.CLK(clknet_leaf_63_clk),
    .D(net1273),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11142_ (.CLK(clknet_leaf_58_clk),
    .D(net1453),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11143_ (.CLK(clknet_leaf_57_clk),
    .D(net2876),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11144_ (.CLK(clknet_leaf_57_clk),
    .D(net2131),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11145_ (.CLK(clknet_leaf_58_clk),
    .D(net305),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11146_ (.CLK(clknet_leaf_58_clk),
    .D(net1140),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11147_ (.CLK(clknet_leaf_59_clk),
    .D(net2463),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11148_ (.CLK(clknet_leaf_56_clk),
    .D(net436),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11149_ (.CLK(clknet_leaf_58_clk),
    .D(net640),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11150_ (.CLK(clknet_leaf_59_clk),
    .D(net2844),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11151_ (.CLK(clknet_leaf_59_clk),
    .D(net2547),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11152_ (.CLK(clknet_leaf_53_clk),
    .D(net917),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11153_ (.CLK(clknet_leaf_53_clk),
    .D(net1083),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11154_ (.CLK(clknet_leaf_49_clk),
    .D(net470),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11155_ (.CLK(clknet_leaf_48_clk),
    .D(net2068),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11156_ (.CLK(clknet_leaf_48_clk),
    .D(net1545),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11157_ (.CLK(clknet_leaf_48_clk),
    .D(net1798),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11158_ (.CLK(clknet_leaf_54_clk),
    .D(net804),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11159_ (.CLK(clknet_leaf_55_clk),
    .D(net193),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11160_ (.CLK(clknet_leaf_55_clk),
    .D(net167),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11161_ (.CLK(clknet_leaf_53_clk),
    .D(net282),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_2 _11162_ (.CLK(clknet_leaf_63_clk),
    .D(net351),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[0] ));
 sky130_fd_sc_hd__dfxtp_2 _11163_ (.CLK(clknet_leaf_64_clk),
    .D(net254),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11164_ (.CLK(clknet_leaf_64_clk),
    .D(net2025),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11165_ (.CLK(clknet_leaf_63_clk),
    .D(net1591),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11166_ (.CLK(clknet_leaf_55_clk),
    .D(net2622),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[4] ));
 sky130_fd_sc_hd__dfxtp_2 _11167_ (.CLK(clknet_leaf_47_clk),
    .D(net2586),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ));
 sky130_fd_sc_hd__dfxtp_2 _11168_ (.CLK(clknet_leaf_47_clk),
    .D(net1053),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11169_ (.CLK(clknet_leaf_44_clk),
    .D(net909),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11170_ (.CLK(clknet_leaf_54_clk),
    .D(net805),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _11171_ (.CLK(clknet_leaf_47_clk),
    .D(net1944),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[9] ));
 sky130_fd_sc_hd__dfxtp_4 _11172_ (.CLK(clknet_leaf_48_clk),
    .D(net944),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ));
 sky130_fd_sc_hd__dfxtp_4 _11173_ (.CLK(clknet_leaf_50_clk),
    .D(net968),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _11174_ (.CLK(clknet_leaf_52_clk),
    .D(net635),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _11175_ (.CLK(clknet_leaf_53_clk),
    .D(net2502),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _11176_ (.CLK(clknet_leaf_52_clk),
    .D(net1745),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[14] ));
 sky130_fd_sc_hd__dfxtp_2 _11177_ (.CLK(clknet_leaf_56_clk),
    .D(net1028),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _11178_ (.CLK(clknet_leaf_56_clk),
    .D(net1055),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[16] ));
 sky130_fd_sc_hd__dfxtp_1 _11179_ (.CLK(clknet_leaf_63_clk),
    .D(net1075),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[17] ));
 sky130_fd_sc_hd__dfxtp_1 _11180_ (.CLK(clknet_leaf_56_clk),
    .D(net965),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[18] ));
 sky130_fd_sc_hd__dfxtp_1 _11181_ (.CLK(clknet_leaf_62_clk),
    .D(net2882),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[19] ));
 sky130_fd_sc_hd__dfxtp_2 _11182_ (.CLK(clknet_leaf_58_clk),
    .D(net1077),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[20] ));
 sky130_fd_sc_hd__dfxtp_2 _11183_ (.CLK(clknet_leaf_57_clk),
    .D(net2062),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[21] ));
 sky130_fd_sc_hd__dfxtp_1 _11184_ (.CLK(clknet_leaf_57_clk),
    .D(net1269),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _11185_ (.CLK(clknet_leaf_59_clk),
    .D(net378),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[23] ));
 sky130_fd_sc_hd__dfxtp_1 _11186_ (.CLK(clknet_leaf_59_clk),
    .D(net400),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[24] ));
 sky130_fd_sc_hd__dfxtp_2 _11187_ (.CLK(clknet_leaf_59_clk),
    .D(net1487),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[25] ));
 sky130_fd_sc_hd__dfxtp_2 _11188_ (.CLK(clknet_leaf_56_clk),
    .D(net1277),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[26] ));
 sky130_fd_sc_hd__dfxtp_1 _11189_ (.CLK(clknet_leaf_58_clk),
    .D(net2122),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[27] ));
 sky130_fd_sc_hd__dfxtp_1 _11190_ (.CLK(clknet_leaf_59_clk),
    .D(net2950),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[28] ));
 sky130_fd_sc_hd__dfxtp_1 _11191_ (.CLK(clknet_leaf_59_clk),
    .D(net2003),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[29] ));
 sky130_fd_sc_hd__dfxtp_2 _11192_ (.CLK(clknet_leaf_57_clk),
    .D(net165),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[30] ));
 sky130_fd_sc_hd__dfxtp_2 _11193_ (.CLK(clknet_leaf_53_clk),
    .D(net847),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[31] ));
 sky130_fd_sc_hd__dfxtp_2 _11194_ (.CLK(clknet_leaf_48_clk),
    .D(net452),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ));
 sky130_fd_sc_hd__dfxtp_2 _11195_ (.CLK(clknet_leaf_48_clk),
    .D(net988),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ));
 sky130_fd_sc_hd__dfxtp_1 _11196_ (.CLK(clknet_leaf_48_clk),
    .D(net2044),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[34] ));
 sky130_fd_sc_hd__dfxtp_4 _11197_ (.CLK(clknet_leaf_48_clk),
    .D(net1033),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ));
 sky130_fd_sc_hd__dfxtp_2 _11198_ (.CLK(clknet_leaf_55_clk),
    .D(net166),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[36] ));
 sky130_fd_sc_hd__dfxtp_1 _11199_ (.CLK(clknet_leaf_55_clk),
    .D(net891),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[37] ));
 sky130_fd_sc_hd__dfxtp_1 _11200_ (.CLK(clknet_leaf_55_clk),
    .D(net880),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[38] ));
 sky130_fd_sc_hd__dfxtp_1 _11201_ (.CLK(clknet_leaf_54_clk),
    .D(net589),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[39] ));
 sky130_fd_sc_hd__dfxtp_2 _11202_ (.CLK(clknet_leaf_51_clk),
    .D(_00030_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _11203_ (.CLK(clknet_leaf_47_clk),
    .D(_00031_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11204_ (.CLK(clknet_leaf_51_clk),
    .D(_00032_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11205_ (.CLK(clknet_leaf_51_clk),
    .D(_00033_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11206_ (.CLK(clknet_leaf_51_clk),
    .D(_00034_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11207_ (.CLK(clknet_leaf_51_clk),
    .D(_00035_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11208_ (.CLK(clknet_leaf_51_clk),
    .D(_00036_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11209_ (.CLK(clknet_leaf_61_clk),
    .D(net3689),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__dfxtp_2 _11210_ (.CLK(clknet_leaf_79_clk),
    .D(net3288),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11211_ (.CLK(clknet_leaf_77_clk),
    .D(net3948),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11212_ (.CLK(clknet_leaf_62_clk),
    .D(net3891),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11213_ (.CLK(clknet_leaf_80_clk),
    .D(net3284),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11214_ (.CLK(clknet_leaf_79_clk),
    .D(net3740),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__dfxtp_2 _11215_ (.CLK(clknet_leaf_79_clk),
    .D(net3828),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__dfxtp_2 _11216_ (.CLK(clknet_leaf_61_clk),
    .D(net3308),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11217_ (.CLK(clknet_leaf_83_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11218_ (.CLK(clknet_leaf_82_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11219_ (.CLK(clknet_leaf_83_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11220_ (.CLK(clknet_leaf_83_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11221_ (.CLK(clknet_leaf_61_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11222_ (.CLK(clknet_leaf_80_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11223_ (.CLK(clknet_leaf_77_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11224_ (.CLK(clknet_leaf_78_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11225_ (.CLK(clknet_leaf_80_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11226_ (.CLK(clknet_leaf_79_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11227_ (.CLK(clknet_leaf_79_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11228_ (.CLK(clknet_leaf_79_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11229_ (.CLK(clknet_leaf_78_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11230_ (.CLK(clknet_leaf_78_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11231_ (.CLK(clknet_leaf_78_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11232_ (.CLK(clknet_leaf_80_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11233_ (.CLK(clknet_leaf_78_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11234_ (.CLK(clknet_leaf_80_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11235_ (.CLK(clknet_leaf_80_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11236_ (.CLK(clknet_leaf_83_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11237_ (.CLK(clknet_leaf_80_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11238_ (.CLK(clknet_leaf_83_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11239_ (.CLK(clknet_leaf_62_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11240_ (.CLK(clknet_leaf_81_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11241_ (.CLK(clknet_leaf_80_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11242_ (.CLK(clknet_leaf_79_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11243_ (.CLK(clknet_leaf_78_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11244_ (.CLK(clknet_leaf_79_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11245_ (.CLK(clknet_leaf_79_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11246_ (.CLK(clknet_leaf_78_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11247_ (.CLK(clknet_leaf_80_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11248_ (.CLK(clknet_leaf_78_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11249_ (.CLK(clknet_leaf_82_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11250_ (.CLK(clknet_leaf_82_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11251_ (.CLK(clknet_leaf_82_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11252_ (.CLK(clknet_leaf_81_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11253_ (.CLK(clknet_leaf_81_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11254_ (.CLK(clknet_leaf_81_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11255_ (.CLK(clknet_leaf_81_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11256_ (.CLK(clknet_leaf_61_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _11257_ (.CLK(clknet_leaf_84_clk),
    .D(net744),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11258_ (.CLK(clknet_leaf_82_clk),
    .D(net2369),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11259_ (.CLK(clknet_leaf_83_clk),
    .D(net2034),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11260_ (.CLK(clknet_leaf_82_clk),
    .D(net670),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11261_ (.CLK(clknet_leaf_61_clk),
    .D(net874),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11262_ (.CLK(clknet_leaf_80_clk),
    .D(net1780),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11263_ (.CLK(clknet_leaf_77_clk),
    .D(net2167),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11264_ (.CLK(clknet_leaf_78_clk),
    .D(net1243),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11265_ (.CLK(clknet_leaf_80_clk),
    .D(net1770),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11266_ (.CLK(clknet_leaf_79_clk),
    .D(net1143),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11267_ (.CLK(clknet_leaf_72_clk),
    .D(net141),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11268_ (.CLK(clknet_leaf_72_clk),
    .D(net130),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11269_ (.CLK(clknet_leaf_78_clk),
    .D(net2728),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11270_ (.CLK(clknet_leaf_78_clk),
    .D(net1284),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11271_ (.CLK(clknet_leaf_78_clk),
    .D(net1600),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11272_ (.CLK(clknet_leaf_62_clk),
    .D(net444),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11273_ (.CLK(clknet_leaf_77_clk),
    .D(net502),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11274_ (.CLK(clknet_leaf_77_clk),
    .D(net531),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11275_ (.CLK(clknet_leaf_83_clk),
    .D(net402),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11276_ (.CLK(clknet_leaf_83_clk),
    .D(net1871),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11277_ (.CLK(clknet_leaf_61_clk),
    .D(net263),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11278_ (.CLK(clknet_leaf_83_clk),
    .D(net1879),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11279_ (.CLK(clknet_leaf_62_clk),
    .D(net1019),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11280_ (.CLK(clknet_leaf_61_clk),
    .D(net186),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11281_ (.CLK(clknet_leaf_80_clk),
    .D(net2431),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11282_ (.CLK(clknet_leaf_79_clk),
    .D(net2911),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11283_ (.CLK(clknet_leaf_78_clk),
    .D(net1271),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11284_ (.CLK(clknet_leaf_79_clk),
    .D(net2303),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11285_ (.CLK(clknet_leaf_79_clk),
    .D(net1901),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11286_ (.CLK(clknet_leaf_78_clk),
    .D(net1767),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11287_ (.CLK(clknet_leaf_78_clk),
    .D(net609),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11288_ (.CLK(clknet_leaf_78_clk),
    .D(net2514),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11289_ (.CLK(clknet_leaf_82_clk),
    .D(net2830),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11290_ (.CLK(clknet_leaf_82_clk),
    .D(net1115),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11291_ (.CLK(clknet_leaf_82_clk),
    .D(net1097),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11292_ (.CLK(clknet_leaf_81_clk),
    .D(net2050),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11293_ (.CLK(clknet_leaf_81_clk),
    .D(net1473),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11294_ (.CLK(clknet_leaf_81_clk),
    .D(net2686),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11295_ (.CLK(clknet_leaf_81_clk),
    .D(net1656),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11296_ (.CLK(clknet_leaf_61_clk),
    .D(net951),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _11297_ (.CLK(clknet_leaf_84_clk),
    .D(net1581),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11298_ (.CLK(clknet_leaf_82_clk),
    .D(net1474),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11299_ (.CLK(clknet_leaf_83_clk),
    .D(net1775),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11300_ (.CLK(clknet_leaf_82_clk),
    .D(net2501),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11301_ (.CLK(clknet_leaf_61_clk),
    .D(net824),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11302_ (.CLK(clknet_leaf_80_clk),
    .D(net2377),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11303_ (.CLK(clknet_leaf_77_clk),
    .D(net2173),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11304_ (.CLK(clknet_leaf_78_clk),
    .D(net1281),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11305_ (.CLK(clknet_leaf_80_clk),
    .D(net2349),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11306_ (.CLK(clknet_leaf_79_clk),
    .D(net1465),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11307_ (.CLK(clknet_leaf_79_clk),
    .D(net539),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11308_ (.CLK(clknet_leaf_73_clk),
    .D(net421),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11309_ (.CLK(clknet_leaf_78_clk),
    .D(net2763),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11310_ (.CLK(clknet_leaf_78_clk),
    .D(net1318),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11311_ (.CLK(clknet_leaf_78_clk),
    .D(net1471),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11312_ (.CLK(clknet_leaf_62_clk),
    .D(net815),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11313_ (.CLK(clknet_leaf_87_clk),
    .D(net517),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11314_ (.CLK(clknet_leaf_77_clk),
    .D(net1168),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11315_ (.CLK(clknet_leaf_87_clk),
    .D(net553),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11316_ (.CLK(clknet_leaf_83_clk),
    .D(net2664),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11317_ (.CLK(clknet_leaf_61_clk),
    .D(net823),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11318_ (.CLK(clknet_leaf_83_clk),
    .D(net1747),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11319_ (.CLK(clknet_leaf_62_clk),
    .D(net813),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11320_ (.CLK(clknet_leaf_81_clk),
    .D(net52),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11321_ (.CLK(clknet_leaf_80_clk),
    .D(net1926),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11322_ (.CLK(clknet_leaf_72_clk),
    .D(net134),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11323_ (.CLK(clknet_leaf_78_clk),
    .D(net1899),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11324_ (.CLK(clknet_leaf_72_clk),
    .D(net140),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11325_ (.CLK(clknet_leaf_79_clk),
    .D(net2326),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11326_ (.CLK(clknet_leaf_78_clk),
    .D(net1278),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11327_ (.CLK(clknet_leaf_78_clk),
    .D(net1653),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11328_ (.CLK(clknet_leaf_77_clk),
    .D(net741),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11329_ (.CLK(clknet_leaf_82_clk),
    .D(net2935),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11330_ (.CLK(clknet_leaf_82_clk),
    .D(net2114),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11331_ (.CLK(clknet_leaf_82_clk),
    .D(net1496),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11332_ (.CLK(clknet_leaf_81_clk),
    .D(net1880),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11333_ (.CLK(clknet_leaf_82_clk),
    .D(net628),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11334_ (.CLK(clknet_leaf_81_clk),
    .D(net1891),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11335_ (.CLK(clknet_leaf_81_clk),
    .D(net1045),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11336_ (.CLK(clknet_leaf_61_clk),
    .D(net912),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_4 _11337_ (.CLK(clknet_leaf_83_clk),
    .D(net311),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ));
 sky130_fd_sc_hd__dfxtp_2 _11338_ (.CLK(clknet_leaf_82_clk),
    .D(net1425),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ));
 sky130_fd_sc_hd__dfxtp_2 _11339_ (.CLK(clknet_leaf_84_clk),
    .D(net540),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11340_ (.CLK(clknet_leaf_83_clk),
    .D(net408),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11341_ (.CLK(clknet_leaf_61_clk),
    .D(net1073),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[4] ));
 sky130_fd_sc_hd__dfxtp_2 _11342_ (.CLK(clknet_leaf_80_clk),
    .D(net1149),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ));
 sky130_fd_sc_hd__dfxtp_2 _11343_ (.CLK(clknet_leaf_87_clk),
    .D(net373),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11344_ (.CLK(clknet_leaf_77_clk),
    .D(net636),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11345_ (.CLK(clknet_leaf_80_clk),
    .D(net2907),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _11346_ (.CLK(clknet_leaf_78_clk),
    .D(net307),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[9] ));
 sky130_fd_sc_hd__dfxtp_2 _11347_ (.CLK(clknet_leaf_79_clk),
    .D(net979),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[10] ));
 sky130_fd_sc_hd__dfxtp_2 _11348_ (.CLK(clknet_leaf_79_clk),
    .D(net328),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _11349_ (.CLK(clknet_leaf_77_clk),
    .D(net611),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _11350_ (.CLK(clknet_leaf_77_clk),
    .D(net616),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _11351_ (.CLK(clknet_leaf_77_clk),
    .D(net627),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[14] ));
 sky130_fd_sc_hd__dfxtp_2 _11352_ (.CLK(clknet_leaf_62_clk),
    .D(net808),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _11353_ (.CLK(clknet_leaf_77_clk),
    .D(net639),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ));
 sky130_fd_sc_hd__dfxtp_2 _11354_ (.CLK(clknet_leaf_87_clk),
    .D(net376),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ));
 sky130_fd_sc_hd__dfxtp_2 _11355_ (.CLK(clknet_leaf_87_clk),
    .D(net1116),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ));
 sky130_fd_sc_hd__dfxtp_1 _11356_ (.CLK(clknet_leaf_83_clk),
    .D(net2742),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[19] ));
 sky130_fd_sc_hd__dfxtp_2 _11357_ (.CLK(clknet_leaf_80_clk),
    .D(net45),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ));
 sky130_fd_sc_hd__dfxtp_2 _11358_ (.CLK(clknet_leaf_87_clk),
    .D(net518),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ));
 sky130_fd_sc_hd__dfxtp_1 _11359_ (.CLK(clknet_leaf_62_clk),
    .D(net802),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _11360_ (.CLK(clknet_leaf_81_clk),
    .D(net2296),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[23] ));
 sky130_fd_sc_hd__dfxtp_1 _11361_ (.CLK(clknet_leaf_80_clk),
    .D(net2917),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[24] ));
 sky130_fd_sc_hd__dfxtp_2 _11362_ (.CLK(clknet_leaf_79_clk),
    .D(net406),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[25] ));
 sky130_fd_sc_hd__dfxtp_2 _11363_ (.CLK(clknet_leaf_77_clk),
    .D(net568),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ));
 sky130_fd_sc_hd__dfxtp_1 _11364_ (.CLK(clknet_leaf_79_clk),
    .D(net542),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[27] ));
 sky130_fd_sc_hd__dfxtp_1 _11365_ (.CLK(clknet_leaf_79_clk),
    .D(net2524),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[28] ));
 sky130_fd_sc_hd__dfxtp_1 _11366_ (.CLK(clknet_leaf_77_clk),
    .D(net637),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[29] ));
 sky130_fd_sc_hd__dfxtp_2 _11367_ (.CLK(clknet_leaf_78_clk),
    .D(net1125),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ));
 sky130_fd_sc_hd__dfxtp_2 _11368_ (.CLK(clknet_leaf_77_clk),
    .D(net1504),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ));
 sky130_fd_sc_hd__dfxtp_2 _11369_ (.CLK(clknet_leaf_82_clk),
    .D(net1106),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ));
 sky130_fd_sc_hd__dfxtp_2 _11370_ (.CLK(clknet_leaf_83_clk),
    .D(net314),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[33] ));
 sky130_fd_sc_hd__dfxtp_1 _11371_ (.CLK(clknet_leaf_82_clk),
    .D(net2187),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[34] ));
 sky130_fd_sc_hd__dfxtp_4 _11372_ (.CLK(clknet_leaf_82_clk),
    .D(net290),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ));
 sky130_fd_sc_hd__dfxtp_2 _11373_ (.CLK(clknet_leaf_81_clk),
    .D(net641),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ));
 sky130_fd_sc_hd__dfxtp_1 _11374_ (.CLK(clknet_leaf_81_clk),
    .D(net1348),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[37] ));
 sky130_fd_sc_hd__dfxtp_1 _11375_ (.CLK(clknet_leaf_80_clk),
    .D(net309),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[38] ));
 sky130_fd_sc_hd__dfxtp_1 _11376_ (.CLK(clknet_leaf_81_clk),
    .D(net53),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[39] ));
 sky130_fd_sc_hd__dfxtp_1 _11377_ (.CLK(clknet_leaf_80_clk),
    .D(_00037_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _11378_ (.CLK(clknet_leaf_83_clk),
    .D(_00038_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11379_ (.CLK(clknet_leaf_83_clk),
    .D(_00039_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11380_ (.CLK(clknet_leaf_83_clk),
    .D(_00040_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11381_ (.CLK(clknet_leaf_83_clk),
    .D(_00041_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11382_ (.CLK(clknet_leaf_80_clk),
    .D(_00042_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11383_ (.CLK(clknet_leaf_80_clk),
    .D(_00043_),
    .Q(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11384_ (.CLK(clknet_leaf_52_clk),
    .D(net3226),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11385_ (.CLK(clknet_leaf_51_clk),
    .D(net3216),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11386_ (.CLK(clknet_leaf_52_clk),
    .D(net3389),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11387_ (.CLK(clknet_leaf_52_clk),
    .D(net3355),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.o[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11388_ (.CLK(clknet_leaf_58_clk),
    .D(net3192),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11389_ (.CLK(clknet_leaf_60_clk),
    .D(net248),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11390_ (.CLK(clknet_leaf_81_clk),
    .D(net3170),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.o[6] ));
 sky130_fd_sc_hd__dfxtp_2 _11391_ (.CLK(clknet_leaf_59_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.o_[7] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11392_ (.CLK(clknet_leaf_52_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11393_ (.CLK(clknet_leaf_52_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11394_ (.CLK(clknet_leaf_51_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11395_ (.CLK(clknet_leaf_51_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11396_ (.CLK(clknet_leaf_49_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11397_ (.CLK(clknet_leaf_48_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11398_ (.CLK(clknet_leaf_50_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11399_ (.CLK(clknet_leaf_48_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11400_ (.CLK(clknet_leaf_50_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11401_ (.CLK(clknet_leaf_50_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11402_ (.CLK(clknet_leaf_50_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11403_ (.CLK(clknet_leaf_49_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11404_ (.CLK(clknet_leaf_49_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11405_ (.CLK(clknet_leaf_49_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11406_ (.CLK(clknet_leaf_49_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11407_ (.CLK(clknet_leaf_49_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11408_ (.CLK(clknet_leaf_57_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11409_ (.CLK(clknet_leaf_57_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11410_ (.CLK(clknet_leaf_57_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11411_ (.CLK(clknet_leaf_58_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11412_ (.CLK(clknet_leaf_60_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11413_ (.CLK(clknet_leaf_60_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11414_ (.CLK(clknet_leaf_60_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11415_ (.CLK(clknet_leaf_60_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11416_ (.CLK(clknet_leaf_83_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11417_ (.CLK(clknet_leaf_82_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11418_ (.CLK(clknet_leaf_82_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11419_ (.CLK(clknet_leaf_81_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11420_ (.CLK(clknet_leaf_58_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11421_ (.CLK(clknet_leaf_58_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11422_ (.CLK(clknet_leaf_60_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11423_ (.CLK(clknet_leaf_59_clk),
    .D(\c.genblk1.genblk1.subs.sw.up.x.selects.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11424_ (.CLK(clknet_leaf_52_clk),
    .D(net1052),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11425_ (.CLK(clknet_leaf_52_clk),
    .D(net1611),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11426_ (.CLK(clknet_leaf_51_clk),
    .D(net2625),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11427_ (.CLK(clknet_leaf_51_clk),
    .D(net2640),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11428_ (.CLK(clknet_leaf_49_clk),
    .D(net2784),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11429_ (.CLK(clknet_leaf_50_clk),
    .D(net623),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11430_ (.CLK(clknet_leaf_50_clk),
    .D(net2385),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11431_ (.CLK(clknet_leaf_49_clk),
    .D(net456),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11432_ (.CLK(clknet_leaf_50_clk),
    .D(net2375),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11433_ (.CLK(clknet_leaf_50_clk),
    .D(net2001),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11434_ (.CLK(clknet_leaf_50_clk),
    .D(net2281),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11435_ (.CLK(clknet_leaf_50_clk),
    .D(net578),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11436_ (.CLK(clknet_leaf_49_clk),
    .D(net2440),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11437_ (.CLK(clknet_leaf_49_clk),
    .D(net2905),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11438_ (.CLK(clknet_leaf_49_clk),
    .D(net1620),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11439_ (.CLK(clknet_leaf_49_clk),
    .D(net1797),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11440_ (.CLK(clknet_leaf_57_clk),
    .D(net1764),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11441_ (.CLK(clknet_leaf_52_clk),
    .D(net100),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11442_ (.CLK(clknet_leaf_58_clk),
    .D(net273),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11443_ (.CLK(clknet_leaf_58_clk),
    .D(net1558),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11444_ (.CLK(clknet_leaf_60_clk),
    .D(net2247),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11445_ (.CLK(clknet_leaf_60_clk),
    .D(net915),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11446_ (.CLK(clknet_leaf_60_clk),
    .D(net994),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11447_ (.CLK(clknet_leaf_60_clk),
    .D(net925),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11448_ (.CLK(clknet_leaf_83_clk),
    .D(net1452),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11449_ (.CLK(clknet_leaf_82_clk),
    .D(net2829),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11450_ (.CLK(clknet_leaf_82_clk),
    .D(net1831),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11451_ (.CLK(clknet_leaf_81_clk),
    .D(net1849),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11452_ (.CLK(clknet_leaf_58_clk),
    .D(net1701),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11453_ (.CLK(clknet_leaf_58_clk),
    .D(net2165),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11454_ (.CLK(clknet_leaf_60_clk),
    .D(net932),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11455_ (.CLK(clknet_leaf_59_clk),
    .D(net1981),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11456_ (.CLK(clknet_leaf_52_clk),
    .D(net1582),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11457_ (.CLK(clknet_leaf_52_clk),
    .D(net1104),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11458_ (.CLK(clknet_leaf_51_clk),
    .D(net1991),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11459_ (.CLK(clknet_leaf_51_clk),
    .D(net1094),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11460_ (.CLK(clknet_leaf_49_clk),
    .D(net2052),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11461_ (.CLK(clknet_leaf_50_clk),
    .D(net1705),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11462_ (.CLK(clknet_leaf_50_clk),
    .D(net2704),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11463_ (.CLK(clknet_leaf_49_clk),
    .D(net2432),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11464_ (.CLK(clknet_leaf_50_clk),
    .D(net2196),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11465_ (.CLK(clknet_leaf_50_clk),
    .D(net1371),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11466_ (.CLK(clknet_leaf_51_clk),
    .D(net572),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11467_ (.CLK(clknet_leaf_50_clk),
    .D(net2470),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11468_ (.CLK(clknet_leaf_49_clk),
    .D(net1820),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11469_ (.CLK(clknet_leaf_49_clk),
    .D(net1706),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11470_ (.CLK(clknet_leaf_50_clk),
    .D(net506),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11471_ (.CLK(clknet_leaf_49_clk),
    .D(net2175),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11472_ (.CLK(clknet_leaf_57_clk),
    .D(net1816),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11473_ (.CLK(clknet_leaf_57_clk),
    .D(net302),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11474_ (.CLK(clknet_leaf_58_clk),
    .D(net2264),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11475_ (.CLK(clknet_leaf_58_clk),
    .D(net2152),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11476_ (.CLK(clknet_leaf_60_clk),
    .D(net1268),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11477_ (.CLK(clknet_leaf_60_clk),
    .D(net882),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11478_ (.CLK(clknet_leaf_60_clk),
    .D(net1461),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11479_ (.CLK(clknet_leaf_60_clk),
    .D(net1241),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11480_ (.CLK(clknet_leaf_83_clk),
    .D(net2866),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11481_ (.CLK(clknet_leaf_82_clk),
    .D(net2029),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11482_ (.CLK(clknet_leaf_84_clk),
    .D(net354),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11483_ (.CLK(clknet_leaf_81_clk),
    .D(net2565),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11484_ (.CLK(clknet_leaf_58_clk),
    .D(net1108),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11485_ (.CLK(clknet_leaf_58_clk),
    .D(net1114),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11486_ (.CLK(clknet_leaf_60_clk),
    .D(net1221),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11487_ (.CLK(clknet_leaf_59_clk),
    .D(net1674),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11488_ (.CLK(clknet_leaf_52_clk),
    .D(net926),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11489_ (.CLK(clknet_leaf_52_clk),
    .D(net936),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11490_ (.CLK(clknet_leaf_52_clk),
    .D(net716),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11491_ (.CLK(clknet_leaf_52_clk),
    .D(net649),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11492_ (.CLK(clknet_leaf_49_clk),
    .D(net1138),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ));
 sky130_fd_sc_hd__dfxtp_2 _11493_ (.CLK(clknet_leaf_50_clk),
    .D(net1127),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11494_ (.CLK(clknet_leaf_51_clk),
    .D(net579),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11495_ (.CLK(clknet_leaf_49_clk),
    .D(net1383),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[7] ));
 sky130_fd_sc_hd__dfxtp_2 _11496_ (.CLK(clknet_leaf_50_clk),
    .D(net1152),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ));
 sky130_fd_sc_hd__dfxtp_2 _11497_ (.CLK(clknet_leaf_51_clk),
    .D(net545),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _11498_ (.CLK(clknet_leaf_51_clk),
    .D(net2800),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _11499_ (.CLK(clknet_leaf_50_clk),
    .D(net1392),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[11] ));
 sky130_fd_sc_hd__dfxtp_2 _11500_ (.CLK(clknet_leaf_49_clk),
    .D(net1986),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ));
 sky130_fd_sc_hd__dfxtp_2 _11501_ (.CLK(clknet_leaf_49_clk),
    .D(net1133),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _11502_ (.CLK(clknet_leaf_50_clk),
    .D(net1917),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _11503_ (.CLK(clknet_leaf_49_clk),
    .D(net1389),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[15] ));
 sky130_fd_sc_hd__dfxtp_1 _11504_ (.CLK(clknet_leaf_57_clk),
    .D(net963),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[16] ));
 sky130_fd_sc_hd__dfxtp_1 _11505_ (.CLK(clknet_leaf_57_clk),
    .D(net1557),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[17] ));
 sky130_fd_sc_hd__dfxtp_1 _11506_ (.CLK(clknet_leaf_58_clk),
    .D(net2388),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[18] ));
 sky130_fd_sc_hd__dfxtp_1 _11507_ (.CLK(clknet_leaf_58_clk),
    .D(net1500),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[19] ));
 sky130_fd_sc_hd__dfxtp_2 _11508_ (.CLK(clknet_leaf_60_clk),
    .D(net1006),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[20] ));
 sky130_fd_sc_hd__dfxtp_1 _11509_ (.CLK(clknet_leaf_60_clk),
    .D(net1821),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[21] ));
 sky130_fd_sc_hd__dfxtp_1 _11510_ (.CLK(clknet_leaf_81_clk),
    .D(net295),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _11511_ (.CLK(clknet_leaf_81_clk),
    .D(net327),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[23] ));
 sky130_fd_sc_hd__dfxtp_2 _11512_ (.CLK(clknet_leaf_84_clk),
    .D(net565),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ));
 sky130_fd_sc_hd__dfxtp_2 _11513_ (.CLK(clknet_leaf_84_clk),
    .D(net403),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ));
 sky130_fd_sc_hd__dfxtp_1 _11514_ (.CLK(clknet_leaf_84_clk),
    .D(net2423),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[26] ));
 sky130_fd_sc_hd__dfxtp_1 _11515_ (.CLK(clknet_leaf_82_clk),
    .D(net446),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[27] ));
 sky130_fd_sc_hd__dfxtp_2 _11516_ (.CLK(clknet_leaf_59_clk),
    .D(net350),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[28] ));
 sky130_fd_sc_hd__dfxtp_1 _11517_ (.CLK(clknet_leaf_58_clk),
    .D(net1704),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[29] ));
 sky130_fd_sc_hd__dfxtp_1 _11518_ (.CLK(clknet_leaf_60_clk),
    .D(net977),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[30] ));
 sky130_fd_sc_hd__dfxtp_1 _11519_ (.CLK(clknet_leaf_60_clk),
    .D(net67),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.o[31] ));
 sky130_fd_sc_hd__dfxtp_4 _11520_ (.CLK(clknet_leaf_61_clk),
    .D(_00044_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _11521_ (.CLK(clknet_leaf_61_clk),
    .D(_00045_),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11522_ (.CLK(clknet_leaf_59_clk),
    .D(net3201),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _11523_ (.CLK(clknet_leaf_59_clk),
    .D(_00047_),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _11524_ (.CLK(clknet_leaf_60_clk),
    .D(net3796),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11525_ (.CLK(clknet_leaf_59_clk),
    .D(_00049_),
    .Q(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11526_ (.CLK(clknet_leaf_49_clk),
    .D(net2971),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _11527_ (.CLK(clknet_leaf_49_clk),
    .D(net2947),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _11528_ (.CLK(clknet_leaf_50_clk),
    .D(net2903),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _11529_ (.CLK(clknet_leaf_51_clk),
    .D(net862),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _11530_ (.CLK(clknet_leaf_92_clk),
    .D(net197),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _11531_ (.CLK(clknet_leaf_93_clk),
    .D(net3107),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _11532_ (.CLK(clknet_leaf_94_clk),
    .D(net2976),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _11533_ (.CLK(clknet_leaf_94_clk),
    .D(net219),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _11534_ (.CLK(clknet_leaf_180_clk),
    .D(net2),
    .Q(\c.cfg_i_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11535_ (.CLK(clknet_leaf_155_clk),
    .D(net3),
    .Q(\c.cfg_i_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11536_ (.CLK(clknet_leaf_154_clk),
    .D(net4),
    .Q(\c.cfg_i_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11537_ (.CLK(clknet_leaf_152_clk),
    .D(net5),
    .Q(\c.cfg_i_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11538_ (.CLK(clknet_leaf_152_clk),
    .D(net6),
    .Q(\c.cfg_i_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11539_ (.CLK(clknet_leaf_189_clk),
    .D(net40),
    .Q(\c.genblk1.genblk1.subs.c0.m[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11540_ (.CLK(clknet_leaf_183_clk),
    .D(net9),
    .Q(\c.genblk1.genblk1.subs.c0.m[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11541_ (.CLK(clknet_leaf_189_clk),
    .D(net38),
    .Q(\c.genblk1.genblk1.subs.c0.grst ));
 sky130_fd_sc_hd__dfxtp_1 _11542_ (.CLK(clknet_leaf_190_clk),
    .D(net10),
    .Q(\c.genblk1.genblk1.subs.c0.rst ));
 sky130_fd_sc_hd__dfxtp_1 _11543_ (.CLK(clknet_leaf_118_clk),
    .D(_00050_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ));
 sky130_fd_sc_hd__dfxtp_1 _11544_ (.CLK(clknet_leaf_85_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11545_ (.CLK(clknet_leaf_85_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11546_ (.CLK(clknet_leaf_85_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11547_ (.CLK(clknet_leaf_85_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11548_ (.CLK(clknet_leaf_91_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11549_ (.CLK(clknet_leaf_85_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11550_ (.CLK(clknet_leaf_91_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11551_ (.CLK(clknet_leaf_85_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11552_ (.CLK(clknet_leaf_83_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11553_ (.CLK(clknet_leaf_83_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11554_ (.CLK(clknet_leaf_86_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11555_ (.CLK(clknet_leaf_86_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11556_ (.CLK(clknet_leaf_84_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11557_ (.CLK(clknet_leaf_84_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11558_ (.CLK(clknet_leaf_84_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11559_ (.CLK(clknet_leaf_85_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11560_ (.CLK(clknet_leaf_90_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11561_ (.CLK(clknet_leaf_90_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11562_ (.CLK(clknet_leaf_90_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11563_ (.CLK(clknet_leaf_86_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11564_ (.CLK(clknet_leaf_92_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11565_ (.CLK(clknet_leaf_91_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11566_ (.CLK(clknet_leaf_92_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11567_ (.CLK(clknet_leaf_91_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11568_ (.CLK(clknet_leaf_89_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11569_ (.CLK(clknet_leaf_89_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11570_ (.CLK(clknet_leaf_86_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11571_ (.CLK(clknet_leaf_90_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11572_ (.CLK(clknet_leaf_93_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11573_ (.CLK(clknet_leaf_93_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11574_ (.CLK(clknet_leaf_94_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11575_ (.CLK(clknet_leaf_93_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11576_ (.CLK(clknet_leaf_76_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11577_ (.CLK(clknet_leaf_73_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11578_ (.CLK(clknet_leaf_77_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11579_ (.CLK(clknet_leaf_76_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11580_ (.CLK(clknet_leaf_77_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11581_ (.CLK(clknet_leaf_87_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11582_ (.CLK(clknet_leaf_76_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11583_ (.CLK(clknet_leaf_87_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _11584_ (.CLK(clknet_leaf_87_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _11585_ (.CLK(clknet_leaf_87_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _11586_ (.CLK(clknet_leaf_86_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _11587_ (.CLK(clknet_leaf_87_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _11588_ (.CLK(clknet_leaf_70_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _11589_ (.CLK(clknet_leaf_70_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _11590_ (.CLK(clknet_leaf_70_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _11591_ (.CLK(clknet_leaf_85_clk),
    .D(net2452),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11592_ (.CLK(clknet_leaf_85_clk),
    .D(net1807),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11593_ (.CLK(clknet_leaf_85_clk),
    .D(net1502),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11594_ (.CLK(clknet_leaf_85_clk),
    .D(net1936),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11595_ (.CLK(clknet_leaf_91_clk),
    .D(net970),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11596_ (.CLK(clknet_leaf_85_clk),
    .D(net1971),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11597_ (.CLK(clknet_leaf_91_clk),
    .D(net985),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11598_ (.CLK(clknet_leaf_91_clk),
    .D(net120),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11599_ (.CLK(clknet_leaf_84_clk),
    .D(net687),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11600_ (.CLK(clknet_leaf_84_clk),
    .D(net560),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11601_ (.CLK(clknet_leaf_86_clk),
    .D(net1025),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11602_ (.CLK(clknet_leaf_86_clk),
    .D(net1027),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11603_ (.CLK(clknet_leaf_84_clk),
    .D(net1800),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11604_ (.CLK(clknet_leaf_84_clk),
    .D(net2607),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11605_ (.CLK(clknet_leaf_84_clk),
    .D(net2793),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11606_ (.CLK(clknet_leaf_84_clk),
    .D(net740),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11607_ (.CLK(clknet_leaf_91_clk),
    .D(net720),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11608_ (.CLK(clknet_leaf_90_clk),
    .D(net2290),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11609_ (.CLK(clknet_leaf_90_clk),
    .D(net1791),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11610_ (.CLK(clknet_leaf_86_clk),
    .D(net933),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11611_ (.CLK(clknet_leaf_92_clk),
    .D(net2766),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11612_ (.CLK(clknet_leaf_91_clk),
    .D(net1099),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11613_ (.CLK(clknet_leaf_92_clk),
    .D(net2058),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11614_ (.CLK(clknet_leaf_91_clk),
    .D(net1062),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11615_ (.CLK(clknet_leaf_89_clk),
    .D(net2279),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11616_ (.CLK(clknet_leaf_92_clk),
    .D(net717),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11617_ (.CLK(clknet_leaf_90_clk),
    .D(net94),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11618_ (.CLK(clknet_leaf_90_clk),
    .D(net1234),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11619_ (.CLK(clknet_leaf_93_clk),
    .D(net1906),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11620_ (.CLK(clknet_leaf_94_clk),
    .D(net371),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11621_ (.CLK(clknet_leaf_94_clk),
    .D(net1177),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11622_ (.CLK(clknet_leaf_93_clk),
    .D(net1294),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11623_ (.CLK(clknet_leaf_76_clk),
    .D(net1081),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11624_ (.CLK(clknet_leaf_75_clk),
    .D(net701),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11625_ (.CLK(clknet_leaf_77_clk),
    .D(net2747),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11626_ (.CLK(clknet_leaf_77_clk),
    .D(net267),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11627_ (.CLK(clknet_leaf_77_clk),
    .D(net1645),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11628_ (.CLK(clknet_leaf_87_clk),
    .D(net2471),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11629_ (.CLK(clknet_leaf_88_clk),
    .D(net91),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11630_ (.CLK(clknet_leaf_87_clk),
    .D(net2718),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _11631_ (.CLK(clknet_leaf_86_clk),
    .D(net800),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _11632_ (.CLK(clknet_leaf_87_clk),
    .D(net1328),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _11633_ (.CLK(clknet_leaf_86_clk),
    .D(net878),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _11634_ (.CLK(clknet_leaf_86_clk),
    .D(net810),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _11635_ (.CLK(clknet_leaf_70_clk),
    .D(net1561),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _11636_ (.CLK(clknet_leaf_70_clk),
    .D(net2636),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _11637_ (.CLK(clknet_leaf_70_clk),
    .D(net1532),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _11638_ (.CLK(clknet_leaf_85_clk),
    .D(net1509),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11639_ (.CLK(clknet_leaf_85_clk),
    .D(net1432),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11640_ (.CLK(clknet_leaf_85_clk),
    .D(net2613),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11641_ (.CLK(clknet_leaf_85_clk),
    .D(net1786),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11642_ (.CLK(clknet_leaf_91_clk),
    .D(net1896),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11643_ (.CLK(clknet_leaf_85_clk),
    .D(net2532),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11644_ (.CLK(clknet_leaf_91_clk),
    .D(net1774),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11645_ (.CLK(clknet_leaf_91_clk),
    .D(net1924),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11646_ (.CLK(clknet_leaf_84_clk),
    .D(net1334),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11647_ (.CLK(clknet_leaf_84_clk),
    .D(net1844),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11648_ (.CLK(clknet_leaf_86_clk),
    .D(net1492),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11649_ (.CLK(clknet_leaf_86_clk),
    .D(net1018),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11650_ (.CLK(clknet_leaf_84_clk),
    .D(net1915),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11651_ (.CLK(clknet_leaf_85_clk),
    .D(net316),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11652_ (.CLK(clknet_leaf_84_clk),
    .D(net2135),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11653_ (.CLK(clknet_leaf_84_clk),
    .D(net1165),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11654_ (.CLK(clknet_leaf_90_clk),
    .D(net324),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11655_ (.CLK(clknet_leaf_90_clk),
    .D(net1610),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11656_ (.CLK(clknet_leaf_90_clk),
    .D(net1447),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11657_ (.CLK(clknet_leaf_86_clk),
    .D(net919),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11658_ (.CLK(clknet_leaf_92_clk),
    .D(net2925),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11659_ (.CLK(clknet_leaf_92_clk),
    .D(net590),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11660_ (.CLK(clknet_leaf_92_clk),
    .D(net2899),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11661_ (.CLK(clknet_leaf_91_clk),
    .D(net961),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11662_ (.CLK(clknet_leaf_92_clk),
    .D(net676),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11663_ (.CLK(clknet_leaf_92_clk),
    .D(net937),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11664_ (.CLK(clknet_leaf_90_clk),
    .D(net1239),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11665_ (.CLK(clknet_leaf_89_clk),
    .D(net398),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11666_ (.CLK(clknet_leaf_94_clk),
    .D(net432),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11667_ (.CLK(clknet_leaf_94_clk),
    .D(net1039),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11668_ (.CLK(clknet_leaf_94_clk),
    .D(net2061),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11669_ (.CLK(clknet_leaf_93_clk),
    .D(net958),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11670_ (.CLK(clknet_leaf_76_clk),
    .D(net904),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11671_ (.CLK(clknet_leaf_75_clk),
    .D(net2518),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11672_ (.CLK(clknet_leaf_77_clk),
    .D(net2339),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11673_ (.CLK(clknet_leaf_76_clk),
    .D(net796),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11674_ (.CLK(clknet_leaf_77_clk),
    .D(net2389),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11675_ (.CLK(clknet_leaf_87_clk),
    .D(net1677),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11676_ (.CLK(clknet_leaf_88_clk),
    .D(net2682),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11677_ (.CLK(clknet_leaf_88_clk),
    .D(net112),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _11678_ (.CLK(clknet_leaf_90_clk),
    .D(net93),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _11679_ (.CLK(clknet_leaf_87_clk),
    .D(net1657),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _11680_ (.CLK(clknet_leaf_90_clk),
    .D(net92),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _11681_ (.CLK(clknet_leaf_87_clk),
    .D(net231),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _11682_ (.CLK(clknet_leaf_70_clk),
    .D(net2840),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _11683_ (.CLK(clknet_leaf_70_clk),
    .D(net2390),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _11684_ (.CLK(clknet_leaf_118_clk),
    .D(net577),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _11685_ (.CLK(clknet_leaf_85_clk),
    .D(net2496),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11686_ (.CLK(clknet_leaf_85_clk),
    .D(net2408),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11687_ (.CLK(clknet_leaf_85_clk),
    .D(net2834),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11688_ (.CLK(clknet_leaf_85_clk),
    .D(net1759),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11689_ (.CLK(clknet_leaf_91_clk),
    .D(net2779),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11690_ (.CLK(clknet_leaf_91_clk),
    .D(net127),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11691_ (.CLK(clknet_leaf_91_clk),
    .D(net2632),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11692_ (.CLK(clknet_leaf_90_clk),
    .D(net346),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11693_ (.CLK(clknet_leaf_84_clk),
    .D(net1520),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _11694_ (.CLK(clknet_leaf_84_clk),
    .D(net1166),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _11695_ (.CLK(clknet_leaf_85_clk),
    .D(net216),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _11696_ (.CLK(clknet_leaf_86_clk),
    .D(net1438),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _11697_ (.CLK(clknet_leaf_84_clk),
    .D(net1760),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _11698_ (.CLK(clknet_leaf_85_clk),
    .D(net2696),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _11699_ (.CLK(clknet_leaf_84_clk),
    .D(net2293),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _11700_ (.CLK(clknet_leaf_85_clk),
    .D(net360),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _11701_ (.CLK(clknet_leaf_90_clk),
    .D(net1067),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11702_ (.CLK(clknet_leaf_90_clk),
    .D(net2703),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11703_ (.CLK(clknet_leaf_89_clk),
    .D(net395),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11704_ (.CLK(clknet_leaf_91_clk),
    .D(net98),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11705_ (.CLK(clknet_leaf_92_clk),
    .D(net1245),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11706_ (.CLK(clknet_leaf_92_clk),
    .D(net2072),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11707_ (.CLK(clknet_leaf_92_clk),
    .D(net2584),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11708_ (.CLK(clknet_leaf_91_clk),
    .D(net1825),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _11709_ (.CLK(clknet_leaf_92_clk),
    .D(net1163),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _11710_ (.CLK(clknet_leaf_93_clk),
    .D(net566),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _11711_ (.CLK(clknet_leaf_90_clk),
    .D(net2085),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _11712_ (.CLK(clknet_leaf_89_clk),
    .D(net2244),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _11713_ (.CLK(clknet_leaf_94_clk),
    .D(net1195),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _11714_ (.CLK(clknet_leaf_94_clk),
    .D(net2023),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _11715_ (.CLK(clknet_leaf_94_clk),
    .D(net2868),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _11716_ (.CLK(clknet_leaf_94_clk),
    .D(net392),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _11717_ (.CLK(clknet_leaf_76_clk),
    .D(net929),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11718_ (.CLK(clknet_leaf_76_clk),
    .D(net321),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11719_ (.CLK(clknet_leaf_77_clk),
    .D(net1988),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11720_ (.CLK(clknet_leaf_76_clk),
    .D(net871),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11721_ (.CLK(clknet_leaf_77_clk),
    .D(net1469),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11722_ (.CLK(clknet_leaf_87_clk),
    .D(net1304),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11723_ (.CLK(clknet_leaf_88_clk),
    .D(net2927),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11724_ (.CLK(clknet_leaf_88_clk),
    .D(net1449),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11725_ (.CLK(clknet_leaf_89_clk),
    .D(net547),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _11726_ (.CLK(clknet_leaf_87_clk),
    .D(net1266),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _11727_ (.CLK(clknet_leaf_90_clk),
    .D(net2617),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _11728_ (.CLK(clknet_leaf_87_clk),
    .D(net2455),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _11729_ (.CLK(clknet_leaf_70_clk),
    .D(net2569),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _11730_ (.CLK(clknet_leaf_70_clk),
    .D(net2360),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _11731_ (.CLK(clknet_leaf_118_clk),
    .D(net2919),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _11732_ (.CLK(clknet_leaf_87_clk),
    .D(_00051_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _11733_ (.CLK(clknet_leaf_87_clk),
    .D(_00052_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11734_ (.CLK(clknet_leaf_87_clk),
    .D(_00053_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11735_ (.CLK(clknet_leaf_86_clk),
    .D(_00054_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11736_ (.CLK(clknet_leaf_86_clk),
    .D(_00055_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11737_ (.CLK(clknet_leaf_86_clk),
    .D(_00056_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _11738_ (.CLK(clknet_leaf_87_clk),
    .D(_00057_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11739_ (.CLK(clknet_leaf_122_clk),
    .D(_00058_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ));
 sky130_fd_sc_hd__dfxtp_1 _11740_ (.CLK(clknet_leaf_71_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11741_ (.CLK(clknet_leaf_71_clk),
    .D(net1822),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11742_ (.CLK(clknet_leaf_71_clk),
    .D(net1575),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11743_ (.CLK(clknet_leaf_70_clk),
    .D(net342),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11744_ (.CLK(clknet_leaf_92_clk),
    .D(_00012_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _11745_ (.CLK(clknet_leaf_92_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11746_ (.CLK(clknet_leaf_93_clk),
    .D(net2986),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11747_ (.CLK(clknet_leaf_93_clk),
    .D(net3043),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11748_ (.CLK(clknet_leaf_92_clk),
    .D(net2993),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11749_ (.CLK(clknet_leaf_87_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11750_ (.CLK(clknet_leaf_93_clk),
    .D(net2983),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11751_ (.CLK(clknet_leaf_93_clk),
    .D(net3089),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11752_ (.CLK(clknet_leaf_93_clk),
    .D(net3088),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11753_ (.CLK(clknet_leaf_88_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _11754_ (.CLK(clknet_leaf_91_clk),
    .D(net3136),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _11755_ (.CLK(clknet_leaf_91_clk),
    .D(net3078),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _11756_ (.CLK(clknet_leaf_91_clk),
    .D(net3063),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _11757_ (.CLK(clknet_leaf_90_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _11758_ (.CLK(clknet_leaf_92_clk),
    .D(net3010),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _11759_ (.CLK(clknet_leaf_92_clk),
    .D(net3087),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _11760_ (.CLK(clknet_leaf_92_clk),
    .D(net3125),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _11761_ (.CLK(clknet_leaf_98_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11762_ (.CLK(clknet_leaf_97_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11763_ (.CLK(clknet_leaf_97_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11764_ (.CLK(clknet_leaf_97_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11765_ (.CLK(clknet_leaf_98_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11766_ (.CLK(clknet_leaf_98_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11767_ (.CLK(clknet_leaf_98_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11768_ (.CLK(clknet_leaf_98_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11769_ (.CLK(clknet_leaf_99_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11770_ (.CLK(clknet_leaf_99_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11771_ (.CLK(clknet_leaf_100_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11772_ (.CLK(clknet_leaf_100_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11773_ (.CLK(clknet_leaf_97_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11774_ (.CLK(clknet_leaf_96_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11775_ (.CLK(clknet_leaf_96_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11776_ (.CLK(clknet_leaf_96_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11777_ (.CLK(clknet_leaf_89_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11778_ (.CLK(clknet_leaf_89_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11779_ (.CLK(clknet_leaf_89_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11780_ (.CLK(clknet_leaf_90_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11781_ (.CLK(clknet_leaf_95_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11782_ (.CLK(clknet_leaf_93_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11783_ (.CLK(clknet_leaf_95_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11784_ (.CLK(clknet_leaf_95_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11785_ (.CLK(clknet_leaf_89_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11786_ (.CLK(clknet_leaf_89_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11787_ (.CLK(clknet_leaf_99_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11788_ (.CLK(clknet_leaf_99_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11789_ (.CLK(clknet_leaf_94_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11790_ (.CLK(clknet_leaf_93_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11791_ (.CLK(clknet_leaf_95_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11792_ (.CLK(clknet_leaf_94_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11793_ (.CLK(clknet_leaf_75_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11794_ (.CLK(clknet_leaf_75_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11795_ (.CLK(clknet_leaf_76_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11796_ (.CLK(clknet_leaf_76_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11797_ (.CLK(clknet_leaf_100_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11798_ (.CLK(clknet_leaf_76_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11799_ (.CLK(clknet_leaf_88_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11800_ (.CLK(clknet_leaf_88_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _11801_ (.CLK(clknet_leaf_88_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _11802_ (.CLK(clknet_leaf_100_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _11803_ (.CLK(clknet_leaf_100_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _11804_ (.CLK(clknet_leaf_100_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _11805_ (.CLK(clknet_leaf_69_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _11806_ (.CLK(clknet_leaf_69_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _11807_ (.CLK(clknet_leaf_69_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _11808_ (.CLK(clknet_leaf_98_clk),
    .D(net2865),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11809_ (.CLK(clknet_leaf_97_clk),
    .D(net2148),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11810_ (.CLK(clknet_leaf_97_clk),
    .D(net1211),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11811_ (.CLK(clknet_leaf_97_clk),
    .D(net1250),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11812_ (.CLK(clknet_leaf_98_clk),
    .D(net2867),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11813_ (.CLK(clknet_leaf_98_clk),
    .D(net2374),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11814_ (.CLK(clknet_leaf_96_clk),
    .D(net333),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11815_ (.CLK(clknet_leaf_98_clk),
    .D(net1491),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11816_ (.CLK(clknet_leaf_99_clk),
    .D(net2552),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11817_ (.CLK(clknet_leaf_99_clk),
    .D(net2550),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11818_ (.CLK(clknet_leaf_99_clk),
    .D(net431),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11819_ (.CLK(clknet_leaf_99_clk),
    .D(net364),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11820_ (.CLK(clknet_leaf_97_clk),
    .D(net2125),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11821_ (.CLK(clknet_leaf_96_clk),
    .D(net1324),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11822_ (.CLK(clknet_leaf_96_clk),
    .D(net2835),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11823_ (.CLK(clknet_leaf_96_clk),
    .D(net2292),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11824_ (.CLK(clknet_leaf_89_clk),
    .D(net2468),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11825_ (.CLK(clknet_leaf_90_clk),
    .D(net529),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11826_ (.CLK(clknet_leaf_89_clk),
    .D(net1965),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11827_ (.CLK(clknet_leaf_89_clk),
    .D(net483),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11828_ (.CLK(clknet_leaf_93_clk),
    .D(net428),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11829_ (.CLK(clknet_leaf_95_clk),
    .D(net404),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11830_ (.CLK(clknet_leaf_94_clk),
    .D(net306),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11831_ (.CLK(clknet_leaf_95_clk),
    .D(net1718),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11832_ (.CLK(clknet_leaf_89_clk),
    .D(net2614),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11833_ (.CLK(clknet_leaf_89_clk),
    .D(net2861),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11834_ (.CLK(clknet_leaf_99_clk),
    .D(net2557),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11835_ (.CLK(clknet_leaf_99_clk),
    .D(net1307),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11836_ (.CLK(clknet_leaf_94_clk),
    .D(net1687),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11837_ (.CLK(clknet_leaf_93_clk),
    .D(net1003),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11838_ (.CLK(clknet_leaf_95_clk),
    .D(net1415),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11839_ (.CLK(clknet_leaf_94_clk),
    .D(net2878),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11840_ (.CLK(clknet_leaf_75_clk),
    .D(net1011),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11841_ (.CLK(clknet_leaf_76_clk),
    .D(net341),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11842_ (.CLK(clknet_leaf_76_clk),
    .D(net2787),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11843_ (.CLK(clknet_leaf_113_clk),
    .D(net101),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11844_ (.CLK(clknet_leaf_101_clk),
    .D(net176),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11845_ (.CLK(clknet_leaf_113_clk),
    .D(net97),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11846_ (.CLK(clknet_leaf_88_clk),
    .D(net2534),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11847_ (.CLK(clknet_leaf_88_clk),
    .D(net2311),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _11848_ (.CLK(clknet_leaf_88_clk),
    .D(net1572),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _11849_ (.CLK(clknet_leaf_100_clk),
    .D(net2141),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _11850_ (.CLK(clknet_leaf_100_clk),
    .D(net1874),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _11851_ (.CLK(clknet_leaf_100_clk),
    .D(net2093),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _11852_ (.CLK(clknet_leaf_69_clk),
    .D(net2420),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _11853_ (.CLK(clknet_leaf_69_clk),
    .D(net2407),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _11854_ (.CLK(clknet_leaf_119_clk),
    .D(net600),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _11855_ (.CLK(clknet_leaf_97_clk),
    .D(net519),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11856_ (.CLK(clknet_leaf_97_clk),
    .D(net2433),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11857_ (.CLK(clknet_leaf_96_clk),
    .D(net613),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11858_ (.CLK(clknet_leaf_97_clk),
    .D(net2254),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11859_ (.CLK(clknet_leaf_98_clk),
    .D(net1619),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11860_ (.CLK(clknet_leaf_98_clk),
    .D(net1569),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11861_ (.CLK(clknet_leaf_96_clk),
    .D(net2393),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11862_ (.CLK(clknet_leaf_98_clk),
    .D(net2757),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11863_ (.CLK(clknet_leaf_99_clk),
    .D(net2426),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11864_ (.CLK(clknet_leaf_99_clk),
    .D(net2874),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11865_ (.CLK(clknet_leaf_99_clk),
    .D(net1285),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11866_ (.CLK(clknet_leaf_99_clk),
    .D(net1574),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11867_ (.CLK(clknet_leaf_97_clk),
    .D(net2288),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11868_ (.CLK(clknet_leaf_96_clk),
    .D(net2822),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11869_ (.CLK(clknet_leaf_96_clk),
    .D(net2409),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11870_ (.CLK(clknet_leaf_96_clk),
    .D(net2382),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11871_ (.CLK(clknet_leaf_89_clk),
    .D(net2765),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11872_ (.CLK(clknet_leaf_90_clk),
    .D(net2233),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11873_ (.CLK(clknet_leaf_89_clk),
    .D(net1710),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11874_ (.CLK(clknet_leaf_90_clk),
    .D(net580),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11875_ (.CLK(clknet_leaf_95_clk),
    .D(net380),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11876_ (.CLK(clknet_leaf_95_clk),
    .D(net898),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11877_ (.CLK(clknet_leaf_95_clk),
    .D(net733),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11878_ (.CLK(clknet_leaf_95_clk),
    .D(net1927),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _11879_ (.CLK(clknet_leaf_89_clk),
    .D(net1593),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11880_ (.CLK(clknet_leaf_99_clk),
    .D(net532),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11881_ (.CLK(clknet_leaf_99_clk),
    .D(net2821),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11882_ (.CLK(clknet_leaf_99_clk),
    .D(net1972),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11883_ (.CLK(clknet_leaf_94_clk),
    .D(net2119),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11884_ (.CLK(clknet_leaf_94_clk),
    .D(net374),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11885_ (.CLK(clknet_leaf_95_clk),
    .D(net1644),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _11886_ (.CLK(clknet_leaf_95_clk),
    .D(net675),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _11887_ (.CLK(clknet_leaf_75_clk),
    .D(net1862),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _11888_ (.CLK(clknet_leaf_75_clk),
    .D(net126),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _11889_ (.CLK(clknet_leaf_76_clk),
    .D(net1410),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _11890_ (.CLK(clknet_leaf_76_clk),
    .D(net292),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _11891_ (.CLK(clknet_leaf_101_clk),
    .D(net2528),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _11892_ (.CLK(clknet_leaf_113_clk),
    .D(net2782),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _11893_ (.CLK(clknet_leaf_88_clk),
    .D(net1694),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _11894_ (.CLK(clknet_leaf_88_clk),
    .D(net2790),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _11895_ (.CLK(clknet_leaf_100_clk),
    .D(net665),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _11896_ (.CLK(clknet_leaf_100_clk),
    .D(net1132),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _11897_ (.CLK(clknet_leaf_100_clk),
    .D(net1110),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _11898_ (.CLK(clknet_leaf_100_clk),
    .D(net1996),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _11899_ (.CLK(clknet_leaf_69_clk),
    .D(net2284),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _11900_ (.CLK(clknet_leaf_69_clk),
    .D(net1748),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _11901_ (.CLK(clknet_leaf_119_clk),
    .D(net1206),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _11902_ (.CLK(clknet_leaf_97_clk),
    .D(net2216),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11903_ (.CLK(clknet_leaf_97_clk),
    .D(net1700),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11904_ (.CLK(clknet_leaf_97_clk),
    .D(net583),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11905_ (.CLK(clknet_leaf_97_clk),
    .D(net2772),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11906_ (.CLK(clknet_leaf_98_clk),
    .D(net1539),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11907_ (.CLK(clknet_leaf_98_clk),
    .D(net2505),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11908_ (.CLK(clknet_leaf_96_clk),
    .D(net2465),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11909_ (.CLK(clknet_leaf_96_clk),
    .D(net417),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11910_ (.CLK(clknet_leaf_99_clk),
    .D(net1885),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _11911_ (.CLK(clknet_leaf_99_clk),
    .D(net2775),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _11912_ (.CLK(clknet_leaf_99_clk),
    .D(net1741),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _11913_ (.CLK(clknet_leaf_99_clk),
    .D(net1288),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _11914_ (.CLK(clknet_leaf_96_clk),
    .D(net673),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _11915_ (.CLK(clknet_leaf_96_clk),
    .D(net2507),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _11916_ (.CLK(clknet_leaf_96_clk),
    .D(net2828),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _11917_ (.CLK(clknet_leaf_96_clk),
    .D(net2859),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _11918_ (.CLK(clknet_leaf_89_clk),
    .D(net1634),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11919_ (.CLK(clknet_leaf_89_clk),
    .D(net410),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11920_ (.CLK(clknet_leaf_89_clk),
    .D(net2574),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11921_ (.CLK(clknet_leaf_90_clk),
    .D(net1559),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11922_ (.CLK(clknet_leaf_95_clk),
    .D(net942),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11923_ (.CLK(clknet_leaf_95_clk),
    .D(net1022),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11924_ (.CLK(clknet_leaf_95_clk),
    .D(net2922),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11925_ (.CLK(clknet_leaf_95_clk),
    .D(net2151),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _11926_ (.CLK(clknet_leaf_99_clk),
    .D(net372),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _11927_ (.CLK(clknet_leaf_99_clk),
    .D(net2294),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _11928_ (.CLK(clknet_leaf_98_clk),
    .D(net681),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _11929_ (.CLK(clknet_leaf_99_clk),
    .D(net2537),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _11930_ (.CLK(clknet_leaf_94_clk),
    .D(net1716),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_2 _11931_ (.CLK(clknet_leaf_94_clk),
    .D(net1049),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _11932_ (.CLK(clknet_leaf_96_clk),
    .D(net329),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _11933_ (.CLK(clknet_leaf_95_clk),
    .D(net1068),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _11934_ (.CLK(clknet_leaf_75_clk),
    .D(net1102),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11935_ (.CLK(clknet_leaf_76_clk),
    .D(net338),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11936_ (.CLK(clknet_leaf_76_clk),
    .D(net2073),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11937_ (.CLK(clknet_leaf_76_clk),
    .D(net927),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11938_ (.CLK(clknet_leaf_100_clk),
    .D(net178),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11939_ (.CLK(clknet_leaf_100_clk),
    .D(net171),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11940_ (.CLK(clknet_leaf_88_clk),
    .D(net2812),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11941_ (.CLK(clknet_leaf_88_clk),
    .D(net2071),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11942_ (.CLK(clknet_leaf_100_clk),
    .D(net2771),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _11943_ (.CLK(clknet_leaf_100_clk),
    .D(net2591),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _11944_ (.CLK(clknet_leaf_100_clk),
    .D(net2099),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _11945_ (.CLK(clknet_leaf_100_clk),
    .D(net2737),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _11946_ (.CLK(clknet_leaf_69_clk),
    .D(net1538),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _11947_ (.CLK(clknet_leaf_69_clk),
    .D(net2370),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _11948_ (.CLK(clknet_leaf_118_clk),
    .D(net476),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _11949_ (.CLK(clknet_leaf_88_clk),
    .D(_00059_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _11950_ (.CLK(clknet_leaf_88_clk),
    .D(_00060_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11951_ (.CLK(clknet_leaf_88_clk),
    .D(_00061_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11952_ (.CLK(clknet_leaf_88_clk),
    .D(_00062_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11953_ (.CLK(clknet_leaf_89_clk),
    .D(_00063_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11954_ (.CLK(clknet_leaf_88_clk),
    .D(_00064_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _11955_ (.CLK(clknet_leaf_88_clk),
    .D(_00065_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11956_ (.CLK(clknet_leaf_70_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11957_ (.CLK(clknet_leaf_70_clk),
    .D(net1808),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11958_ (.CLK(clknet_leaf_70_clk),
    .D(net1407),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11959_ (.CLK(clknet_leaf_70_clk),
    .D(net1755),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11960_ (.CLK(clknet_leaf_100_clk),
    .D(_00013_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _11961_ (.CLK(clknet_leaf_99_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11962_ (.CLK(clknet_leaf_96_clk),
    .D(net2989),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11963_ (.CLK(clknet_leaf_96_clk),
    .D(net3074),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11964_ (.CLK(clknet_leaf_96_clk),
    .D(net3103),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11965_ (.CLK(clknet_leaf_88_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11966_ (.CLK(clknet_leaf_93_clk),
    .D(net3144),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11967_ (.CLK(clknet_leaf_95_clk),
    .D(net2968),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _11968_ (.CLK(clknet_leaf_95_clk),
    .D(net3026),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _11969_ (.CLK(clknet_leaf_88_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _11970_ (.CLK(clknet_leaf_89_clk),
    .D(net3106),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _11971_ (.CLK(clknet_leaf_93_clk),
    .D(net3002),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _11972_ (.CLK(clknet_leaf_93_clk),
    .D(net3049),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _11973_ (.CLK(clknet_leaf_98_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _11974_ (.CLK(clknet_leaf_96_clk),
    .D(net2998),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _11975_ (.CLK(clknet_leaf_96_clk),
    .D(net3105),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _11976_ (.CLK(clknet_leaf_96_clk),
    .D(net3102),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _11977_ (.CLK(clknet_leaf_98_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11978_ (.CLK(clknet_leaf_98_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11979_ (.CLK(clknet_leaf_97_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11980_ (.CLK(clknet_leaf_97_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11981_ (.CLK(clknet_leaf_103_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11982_ (.CLK(clknet_leaf_103_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11983_ (.CLK(clknet_leaf_103_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11984_ (.CLK(clknet_leaf_103_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11985_ (.CLK(clknet_leaf_113_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11986_ (.CLK(clknet_leaf_113_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11987_ (.CLK(clknet_leaf_113_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11988_ (.CLK(clknet_leaf_101_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11989_ (.CLK(clknet_leaf_101_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11990_ (.CLK(clknet_leaf_100_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11991_ (.CLK(clknet_leaf_98_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11992_ (.CLK(clknet_leaf_101_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11993_ (.CLK(clknet_leaf_112_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11994_ (.CLK(clknet_leaf_112_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11995_ (.CLK(clknet_leaf_112_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11996_ (.CLK(clknet_leaf_101_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11997_ (.CLK(clknet_leaf_104_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11998_ (.CLK(clknet_leaf_104_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11999_ (.CLK(clknet_leaf_104_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12000_ (.CLK(clknet_leaf_103_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12001_ (.CLK(clknet_leaf_112_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12002_ (.CLK(clknet_leaf_112_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12003_ (.CLK(clknet_leaf_113_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12004_ (.CLK(clknet_leaf_101_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12005_ (.CLK(clknet_leaf_104_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12006_ (.CLK(clknet_leaf_104_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12007_ (.CLK(clknet_leaf_105_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12008_ (.CLK(clknet_leaf_104_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12009_ (.CLK(clknet_leaf_75_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12010_ (.CLK(clknet_leaf_75_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12011_ (.CLK(clknet_leaf_75_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12012_ (.CLK(clknet_leaf_114_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12013_ (.CLK(clknet_leaf_74_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12014_ (.CLK(clknet_leaf_114_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12015_ (.CLK(clknet_leaf_115_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12016_ (.CLK(clknet_leaf_114_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12017_ (.CLK(clknet_leaf_113_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12018_ (.CLK(clknet_leaf_113_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12019_ (.CLK(clknet_leaf_74_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12020_ (.CLK(clknet_leaf_113_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12021_ (.CLK(clknet_leaf_70_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12022_ (.CLK(clknet_leaf_118_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12023_ (.CLK(clknet_leaf_118_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12024_ (.CLK(clknet_leaf_98_clk),
    .D(net2301),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12025_ (.CLK(clknet_leaf_97_clk),
    .D(net361),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12026_ (.CLK(clknet_leaf_97_clk),
    .D(net1664),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12027_ (.CLK(clknet_leaf_103_clk),
    .D(net232),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12028_ (.CLK(clknet_leaf_102_clk),
    .D(net272),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12029_ (.CLK(clknet_leaf_103_clk),
    .D(net1367),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12030_ (.CLK(clknet_leaf_103_clk),
    .D(net1091),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12031_ (.CLK(clknet_leaf_103_clk),
    .D(net1041),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12032_ (.CLK(clknet_leaf_101_clk),
    .D(net621),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12033_ (.CLK(clknet_leaf_101_clk),
    .D(net496),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12034_ (.CLK(clknet_leaf_113_clk),
    .D(net1345),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12035_ (.CLK(clknet_leaf_101_clk),
    .D(net2523),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12036_ (.CLK(clknet_leaf_101_clk),
    .D(net2914),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12037_ (.CLK(clknet_leaf_100_clk),
    .D(net2581),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12038_ (.CLK(clknet_leaf_98_clk),
    .D(net2579),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12039_ (.CLK(clknet_leaf_102_clk),
    .D(net552),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12040_ (.CLK(clknet_leaf_112_clk),
    .D(net1643),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12041_ (.CLK(clknet_leaf_102_clk),
    .D(net281),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12042_ (.CLK(clknet_leaf_112_clk),
    .D(net1691),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12043_ (.CLK(clknet_leaf_101_clk),
    .D(net1796),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12044_ (.CLK(clknet_leaf_104_clk),
    .D(net1932),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12045_ (.CLK(clknet_leaf_104_clk),
    .D(net1563),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12046_ (.CLK(clknet_leaf_104_clk),
    .D(net1267),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12047_ (.CLK(clknet_leaf_104_clk),
    .D(net237),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12048_ (.CLK(clknet_leaf_112_clk),
    .D(net1612),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12049_ (.CLK(clknet_leaf_112_clk),
    .D(net1578),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12050_ (.CLK(clknet_leaf_113_clk),
    .D(net1983),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12051_ (.CLK(clknet_leaf_101_clk),
    .D(net2416),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12052_ (.CLK(clknet_leaf_104_clk),
    .D(net1421),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12053_ (.CLK(clknet_leaf_106_clk),
    .D(net447),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12054_ (.CLK(clknet_leaf_105_clk),
    .D(net1765),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12055_ (.CLK(clknet_leaf_105_clk),
    .D(net399),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12056_ (.CLK(clknet_leaf_75_clk),
    .D(net1069),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12057_ (.CLK(clknet_leaf_75_clk),
    .D(net1338),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12058_ (.CLK(clknet_leaf_74_clk),
    .D(net357),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12059_ (.CLK(clknet_leaf_114_clk),
    .D(net1226),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12060_ (.CLK(clknet_leaf_114_clk),
    .D(net705),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12061_ (.CLK(clknet_leaf_114_clk),
    .D(net939),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12062_ (.CLK(clknet_leaf_115_clk),
    .D(net1743),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12063_ (.CLK(clknet_leaf_114_clk),
    .D(net1089),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12064_ (.CLK(clknet_leaf_114_clk),
    .D(net173),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12065_ (.CLK(clknet_leaf_113_clk),
    .D(net2558),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12066_ (.CLK(clknet_leaf_74_clk),
    .D(net1161),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12067_ (.CLK(clknet_leaf_113_clk),
    .D(net2684),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12068_ (.CLK(clknet_leaf_70_clk),
    .D(net2396),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12069_ (.CLK(clknet_leaf_118_clk),
    .D(net1731),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12070_ (.CLK(clknet_leaf_118_clk),
    .D(net1424),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12071_ (.CLK(clknet_leaf_98_clk),
    .D(net2643),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12072_ (.CLK(clknet_leaf_97_clk),
    .D(net1189),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12073_ (.CLK(clknet_leaf_103_clk),
    .D(net255),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12074_ (.CLK(clknet_leaf_97_clk),
    .D(net153),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12075_ (.CLK(clknet_leaf_103_clk),
    .D(net793),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12076_ (.CLK(clknet_leaf_103_clk),
    .D(net1886),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12077_ (.CLK(clknet_leaf_103_clk),
    .D(net893),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12078_ (.CLK(clknet_leaf_103_clk),
    .D(net883),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12079_ (.CLK(clknet_leaf_101_clk),
    .D(net2429),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12080_ (.CLK(clknet_leaf_101_clk),
    .D(net2676),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12081_ (.CLK(clknet_leaf_113_clk),
    .D(net1354),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12082_ (.CLK(clknet_leaf_101_clk),
    .D(net2714),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12083_ (.CLK(clknet_leaf_100_clk),
    .D(net180),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12084_ (.CLK(clknet_leaf_101_clk),
    .D(net185),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12085_ (.CLK(clknet_leaf_98_clk),
    .D(net1689),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12086_ (.CLK(clknet_leaf_102_clk),
    .D(net1830),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12087_ (.CLK(clknet_leaf_112_clk),
    .D(net934),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12088_ (.CLK(clknet_leaf_102_clk),
    .D(net1959),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12089_ (.CLK(clknet_leaf_102_clk),
    .D(net262),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12090_ (.CLK(clknet_leaf_102_clk),
    .D(net574),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12091_ (.CLK(clknet_leaf_104_clk),
    .D(net2934),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12092_ (.CLK(clknet_leaf_104_clk),
    .D(net1289),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12093_ (.CLK(clknet_leaf_104_clk),
    .D(net1864),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12094_ (.CLK(clknet_leaf_104_clk),
    .D(net1282),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12095_ (.CLK(clknet_leaf_112_clk),
    .D(net1175),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12096_ (.CLK(clknet_leaf_102_clk),
    .D(net388),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12097_ (.CLK(clknet_leaf_113_clk),
    .D(net1340),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12098_ (.CLK(clknet_leaf_101_clk),
    .D(net1399),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12099_ (.CLK(clknet_leaf_104_clk),
    .D(net1749),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12100_ (.CLK(clknet_leaf_106_clk),
    .D(net2918),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12101_ (.CLK(clknet_leaf_105_clk),
    .D(net2434),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12102_ (.CLK(clknet_leaf_104_clk),
    .D(net525),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12103_ (.CLK(clknet_leaf_75_clk),
    .D(net2743),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12104_ (.CLK(clknet_leaf_75_clk),
    .D(net2660),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12105_ (.CLK(clknet_leaf_74_clk),
    .D(net1688),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12106_ (.CLK(clknet_leaf_114_clk),
    .D(net1497),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12107_ (.CLK(clknet_leaf_114_clk),
    .D(net1723),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12108_ (.CLK(clknet_leaf_114_clk),
    .D(net955),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12109_ (.CLK(clknet_leaf_114_clk),
    .D(net783),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12110_ (.CLK(clknet_leaf_114_clk),
    .D(net2097),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12111_ (.CLK(clknet_leaf_113_clk),
    .D(net121),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12112_ (.CLK(clknet_leaf_113_clk),
    .D(net1872),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12113_ (.CLK(clknet_leaf_75_clk),
    .D(net664),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12114_ (.CLK(clknet_leaf_113_clk),
    .D(net2193),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12115_ (.CLK(clknet_leaf_70_clk),
    .D(net2327),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12116_ (.CLK(clknet_leaf_118_clk),
    .D(net1990),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12117_ (.CLK(clknet_leaf_118_clk),
    .D(net2230),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12118_ (.CLK(clknet_leaf_98_clk),
    .D(net1188),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12119_ (.CLK(clknet_leaf_97_clk),
    .D(net2734),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12120_ (.CLK(clknet_leaf_97_clk),
    .D(net162),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12121_ (.CLK(clknet_leaf_97_clk),
    .D(net1566),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12122_ (.CLK(clknet_leaf_103_clk),
    .D(net1601),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12123_ (.CLK(clknet_leaf_103_clk),
    .D(net1632),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12124_ (.CLK(clknet_leaf_103_clk),
    .D(net2443),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12125_ (.CLK(clknet_leaf_103_clk),
    .D(net2123),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12126_ (.CLK(clknet_leaf_101_clk),
    .D(net2906),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12127_ (.CLK(clknet_leaf_101_clk),
    .D(net1935),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12128_ (.CLK(clknet_leaf_100_clk),
    .D(net175),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12129_ (.CLK(clknet_leaf_101_clk),
    .D(net2491),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12130_ (.CLK(clknet_leaf_101_clk),
    .D(net177),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12131_ (.CLK(clknet_leaf_101_clk),
    .D(net1240),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12132_ (.CLK(clknet_leaf_98_clk),
    .D(net2593),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12133_ (.CLK(clknet_leaf_103_clk),
    .D(net782),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _12134_ (.CLK(clknet_leaf_102_clk),
    .D(net264),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12135_ (.CLK(clknet_leaf_102_clk),
    .D(net1440),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12136_ (.CLK(clknet_leaf_102_clk),
    .D(net1974),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12137_ (.CLK(clknet_leaf_102_clk),
    .D(net1964),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _12138_ (.CLK(clknet_leaf_104_clk),
    .D(net2666),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12139_ (.CLK(clknet_leaf_104_clk),
    .D(net2871),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12140_ (.CLK(clknet_leaf_104_clk),
    .D(net2937),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12141_ (.CLK(clknet_leaf_104_clk),
    .D(net2435),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12142_ (.CLK(clknet_leaf_112_clk),
    .D(net1515),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12143_ (.CLK(clknet_leaf_102_clk),
    .D(net2166),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12144_ (.CLK(clknet_leaf_113_clk),
    .D(net1480),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12145_ (.CLK(clknet_leaf_101_clk),
    .D(net1909),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12146_ (.CLK(clknet_leaf_104_clk),
    .D(net1436),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_2 _12147_ (.CLK(clknet_leaf_104_clk),
    .D(net638),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12148_ (.CLK(clknet_leaf_104_clk),
    .D(net592),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12149_ (.CLK(clknet_leaf_104_clk),
    .D(net2953),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12150_ (.CLK(clknet_leaf_75_clk),
    .D(net2391),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12151_ (.CLK(clknet_leaf_75_clk),
    .D(net1131),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12152_ (.CLK(clknet_leaf_75_clk),
    .D(net729),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12153_ (.CLK(clknet_leaf_114_clk),
    .D(net947),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12154_ (.CLK(clknet_leaf_114_clk),
    .D(net940),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12155_ (.CLK(clknet_leaf_115_clk),
    .D(net298),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12156_ (.CLK(clknet_leaf_114_clk),
    .D(net1665),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12157_ (.CLK(clknet_leaf_113_clk),
    .D(net142),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12158_ (.CLK(clknet_leaf_113_clk),
    .D(net1404),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12159_ (.CLK(clknet_leaf_113_clk),
    .D(net2877),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12160_ (.CLK(clknet_leaf_113_clk),
    .D(net131),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12161_ (.CLK(clknet_leaf_113_clk),
    .D(net1525),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12162_ (.CLK(clknet_leaf_70_clk),
    .D(net1884),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _12163_ (.CLK(clknet_leaf_118_clk),
    .D(net2442),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _12164_ (.CLK(clknet_leaf_118_clk),
    .D(net2817),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _12165_ (.CLK(clknet_leaf_115_clk),
    .D(_00066_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _12166_ (.CLK(clknet_leaf_114_clk),
    .D(_00067_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12167_ (.CLK(clknet_leaf_114_clk),
    .D(_00068_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12168_ (.CLK(clknet_leaf_114_clk),
    .D(_00069_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12169_ (.CLK(clknet_leaf_112_clk),
    .D(_00070_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12170_ (.CLK(clknet_leaf_112_clk),
    .D(_00071_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12171_ (.CLK(clknet_leaf_112_clk),
    .D(_00072_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12172_ (.CLK(clknet_leaf_74_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12173_ (.CLK(clknet_leaf_70_clk),
    .D(net397),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12174_ (.CLK(clknet_leaf_115_clk),
    .D(net549),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12175_ (.CLK(clknet_leaf_115_clk),
    .D(net1818),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12176_ (.CLK(clknet_leaf_102_clk),
    .D(_00014_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _12177_ (.CLK(clknet_leaf_102_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12178_ (.CLK(clknet_leaf_102_clk),
    .D(net3085),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12179_ (.CLK(clknet_leaf_102_clk),
    .D(net3059),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12180_ (.CLK(clknet_leaf_102_clk),
    .D(net3050),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12181_ (.CLK(clknet_leaf_114_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12182_ (.CLK(clknet_leaf_102_clk),
    .D(net2960),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12183_ (.CLK(clknet_leaf_105_clk),
    .D(net2978),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12184_ (.CLK(clknet_leaf_102_clk),
    .D(net2994),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12185_ (.CLK(clknet_leaf_114_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12186_ (.CLK(clknet_leaf_102_clk),
    .D(net2954),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12187_ (.CLK(clknet_leaf_105_clk),
    .D(net2981),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12188_ (.CLK(clknet_leaf_102_clk),
    .D(net2984),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12189_ (.CLK(clknet_leaf_101_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12190_ (.CLK(clknet_leaf_102_clk),
    .D(net3007),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12191_ (.CLK(clknet_leaf_103_clk),
    .D(net3082),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12192_ (.CLK(clknet_leaf_105_clk),
    .D(net2973),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12193_ (.CLK(clknet_leaf_106_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12194_ (.CLK(clknet_leaf_108_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12195_ (.CLK(clknet_leaf_106_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12196_ (.CLK(clknet_leaf_106_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12197_ (.CLK(clknet_leaf_106_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12198_ (.CLK(clknet_leaf_108_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12199_ (.CLK(clknet_leaf_108_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12200_ (.CLK(clknet_leaf_106_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12201_ (.CLK(clknet_leaf_116_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12202_ (.CLK(clknet_leaf_116_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12203_ (.CLK(clknet_leaf_110_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12204_ (.CLK(clknet_leaf_116_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12205_ (.CLK(clknet_leaf_107_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12206_ (.CLK(clknet_leaf_107_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12207_ (.CLK(clknet_leaf_107_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12208_ (.CLK(clknet_leaf_107_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12209_ (.CLK(clknet_leaf_110_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12210_ (.CLK(clknet_leaf_110_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12211_ (.CLK(clknet_leaf_109_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12212_ (.CLK(clknet_leaf_110_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12213_ (.CLK(clknet_leaf_105_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12214_ (.CLK(clknet_leaf_105_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12215_ (.CLK(clknet_leaf_105_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12216_ (.CLK(clknet_leaf_105_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12217_ (.CLK(clknet_leaf_110_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12218_ (.CLK(clknet_leaf_110_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12219_ (.CLK(clknet_leaf_109_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12220_ (.CLK(clknet_leaf_110_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12221_ (.CLK(clknet_leaf_111_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12222_ (.CLK(clknet_leaf_112_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12223_ (.CLK(clknet_leaf_111_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12224_ (.CLK(clknet_leaf_111_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12225_ (.CLK(clknet_leaf_74_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12226_ (.CLK(clknet_leaf_74_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12227_ (.CLK(clknet_leaf_74_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12228_ (.CLK(clknet_leaf_115_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12229_ (.CLK(clknet_leaf_115_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12230_ (.CLK(clknet_leaf_115_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12231_ (.CLK(clknet_leaf_115_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12232_ (.CLK(clknet_leaf_117_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12233_ (.CLK(clknet_leaf_117_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12234_ (.CLK(clknet_leaf_117_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12235_ (.CLK(clknet_leaf_117_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12236_ (.CLK(clknet_leaf_116_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12237_ (.CLK(clknet_leaf_119_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12238_ (.CLK(clknet_leaf_119_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12239_ (.CLK(clknet_leaf_118_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12240_ (.CLK(clknet_leaf_106_clk),
    .D(net2497),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12241_ (.CLK(clknet_leaf_105_clk),
    .D(net179),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12242_ (.CLK(clknet_leaf_106_clk),
    .D(net2931),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12243_ (.CLK(clknet_leaf_106_clk),
    .D(net1433),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12244_ (.CLK(clknet_leaf_106_clk),
    .D(net1788),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12245_ (.CLK(clknet_leaf_107_clk),
    .D(net214),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12246_ (.CLK(clknet_leaf_107_clk),
    .D(net199),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12247_ (.CLK(clknet_leaf_106_clk),
    .D(net2685),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12248_ (.CLK(clknet_leaf_116_clk),
    .D(net1840),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12249_ (.CLK(clknet_leaf_116_clk),
    .D(net1042),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12250_ (.CLK(clknet_leaf_110_clk),
    .D(net1720),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12251_ (.CLK(clknet_leaf_110_clk),
    .D(net139),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12252_ (.CLK(clknet_leaf_107_clk),
    .D(net2228),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12253_ (.CLK(clknet_leaf_107_clk),
    .D(net2234),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12254_ (.CLK(clknet_leaf_107_clk),
    .D(net2540),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12255_ (.CLK(clknet_leaf_107_clk),
    .D(net1861),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12256_ (.CLK(clknet_leaf_109_clk),
    .D(net795),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12257_ (.CLK(clknet_leaf_109_clk),
    .D(net784),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12258_ (.CLK(clknet_leaf_109_clk),
    .D(net1293),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12259_ (.CLK(clknet_leaf_110_clk),
    .D(net1490),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12260_ (.CLK(clknet_leaf_105_clk),
    .D(net2106),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12261_ (.CLK(clknet_leaf_105_clk),
    .D(net2266),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12262_ (.CLK(clknet_leaf_106_clk),
    .D(net415),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12263_ (.CLK(clknet_leaf_105_clk),
    .D(net1486),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12264_ (.CLK(clknet_leaf_110_clk),
    .D(net1295),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12265_ (.CLK(clknet_leaf_111_clk),
    .D(net702),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12266_ (.CLK(clknet_leaf_109_clk),
    .D(net1516),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12267_ (.CLK(clknet_leaf_110_clk),
    .D(net1588),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12268_ (.CLK(clknet_leaf_112_clk),
    .D(net454),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12269_ (.CLK(clknet_leaf_111_clk),
    .D(net379),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12270_ (.CLK(clknet_leaf_111_clk),
    .D(net953),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12271_ (.CLK(clknet_leaf_111_clk),
    .D(net1484),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12272_ (.CLK(clknet_leaf_74_clk),
    .D(net2939),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12273_ (.CLK(clknet_leaf_74_clk),
    .D(net1182),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12274_ (.CLK(clknet_leaf_74_clk),
    .D(net2004),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12275_ (.CLK(clknet_leaf_115_clk),
    .D(net1692),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12276_ (.CLK(clknet_leaf_115_clk),
    .D(net1351),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12277_ (.CLK(clknet_leaf_115_clk),
    .D(net2811),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12278_ (.CLK(clknet_leaf_115_clk),
    .D(net2576),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12279_ (.CLK(clknet_leaf_117_clk),
    .D(net1835),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12280_ (.CLK(clknet_leaf_118_clk),
    .D(net728),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12281_ (.CLK(clknet_leaf_116_clk),
    .D(net776),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12282_ (.CLK(clknet_leaf_117_clk),
    .D(net2712),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12283_ (.CLK(clknet_leaf_116_clk),
    .D(net1420),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12284_ (.CLK(clknet_leaf_119_clk),
    .D(net1696),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12285_ (.CLK(clknet_leaf_118_clk),
    .D(net625),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12286_ (.CLK(clknet_leaf_118_clk),
    .D(net1485),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12287_ (.CLK(clknet_leaf_106_clk),
    .D(net2791),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12288_ (.CLK(clknet_leaf_105_clk),
    .D(net2522),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12289_ (.CLK(clknet_leaf_106_clk),
    .D(net2608),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12290_ (.CLK(clknet_leaf_106_clk),
    .D(net2898),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12291_ (.CLK(clknet_leaf_106_clk),
    .D(net1427),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12292_ (.CLK(clknet_leaf_108_clk),
    .D(net997),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12293_ (.CLK(clknet_leaf_107_clk),
    .D(net2164),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12294_ (.CLK(clknet_leaf_106_clk),
    .D(net1426),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12295_ (.CLK(clknet_leaf_110_clk),
    .D(net133),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12296_ (.CLK(clknet_leaf_116_clk),
    .D(net1103),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12297_ (.CLK(clknet_leaf_110_clk),
    .D(net2631),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12298_ (.CLK(clknet_leaf_116_clk),
    .D(net163),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12299_ (.CLK(clknet_leaf_107_clk),
    .D(net1503),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12300_ (.CLK(clknet_leaf_107_clk),
    .D(net2735),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12301_ (.CLK(clknet_leaf_107_clk),
    .D(net1130),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12302_ (.CLK(clknet_leaf_107_clk),
    .D(net1129),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12303_ (.CLK(clknet_leaf_109_clk),
    .D(net896),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12304_ (.CLK(clknet_leaf_109_clk),
    .D(net875),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12305_ (.CLK(clknet_leaf_109_clk),
    .D(net854),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12306_ (.CLK(clknet_leaf_110_clk),
    .D(net1973),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12307_ (.CLK(clknet_leaf_105_clk),
    .D(net2909),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12308_ (.CLK(clknet_leaf_105_clk),
    .D(net1768),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12309_ (.CLK(clknet_leaf_106_clk),
    .D(net1417),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12310_ (.CLK(clknet_leaf_105_clk),
    .D(net2769),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12311_ (.CLK(clknet_leaf_110_clk),
    .D(net1185),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12312_ (.CLK(clknet_leaf_111_clk),
    .D(net952),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12313_ (.CLK(clknet_leaf_109_clk),
    .D(net1044),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12314_ (.CLK(clknet_leaf_110_clk),
    .D(net2555),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12315_ (.CLK(clknet_leaf_112_clk),
    .D(net938),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12316_ (.CLK(clknet_leaf_112_clk),
    .D(net682),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12317_ (.CLK(clknet_leaf_111_clk),
    .D(net1510),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12318_ (.CLK(clknet_leaf_112_clk),
    .D(net538),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12319_ (.CLK(clknet_leaf_74_clk),
    .D(net1792),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12320_ (.CLK(clknet_leaf_74_clk),
    .D(net2302),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12321_ (.CLK(clknet_leaf_74_clk),
    .D(net1622),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12322_ (.CLK(clknet_leaf_115_clk),
    .D(net2113),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12323_ (.CLK(clknet_leaf_115_clk),
    .D(net2554),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12324_ (.CLK(clknet_leaf_115_clk),
    .D(net2019),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12325_ (.CLK(clknet_leaf_115_clk),
    .D(net2606),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12326_ (.CLK(clknet_leaf_118_clk),
    .D(net697),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12327_ (.CLK(clknet_leaf_117_clk),
    .D(net458),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12328_ (.CLK(clknet_leaf_117_clk),
    .D(net253),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12329_ (.CLK(clknet_leaf_117_clk),
    .D(net2321),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12330_ (.CLK(clknet_leaf_116_clk),
    .D(net996),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12331_ (.CLK(clknet_leaf_119_clk),
    .D(net1346),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12332_ (.CLK(clknet_leaf_118_clk),
    .D(net2055),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12333_ (.CLK(clknet_leaf_118_clk),
    .D(net1229),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12334_ (.CLK(clknet_leaf_106_clk),
    .D(net2894),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12335_ (.CLK(clknet_leaf_106_clk),
    .D(net575),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12336_ (.CLK(clknet_leaf_106_clk),
    .D(net2921),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12337_ (.CLK(clknet_leaf_106_clk),
    .D(net2896),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12338_ (.CLK(clknet_leaf_107_clk),
    .D(net674),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12339_ (.CLK(clknet_leaf_108_clk),
    .D(net873),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12340_ (.CLK(clknet_leaf_108_clk),
    .D(net1156),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12341_ (.CLK(clknet_leaf_106_clk),
    .D(net2202),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12342_ (.CLK(clknet_leaf_110_clk),
    .D(net1385),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12343_ (.CLK(clknet_leaf_116_clk),
    .D(net908),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12344_ (.CLK(clknet_leaf_110_clk),
    .D(net1995),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12345_ (.CLK(clknet_leaf_110_clk),
    .D(net137),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12346_ (.CLK(clknet_leaf_107_clk),
    .D(net2018),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12347_ (.CLK(clknet_leaf_107_clk),
    .D(net2304),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12348_ (.CLK(clknet_leaf_107_clk),
    .D(net1550),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12349_ (.CLK(clknet_leaf_107_clk),
    .D(net1329),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _12350_ (.CLK(clknet_leaf_108_clk),
    .D(net567),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12351_ (.CLK(clknet_leaf_109_clk),
    .D(net876),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12352_ (.CLK(clknet_leaf_108_clk),
    .D(net698),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12353_ (.CLK(clknet_leaf_110_clk),
    .D(net1209),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _12354_ (.CLK(clknet_leaf_105_clk),
    .D(net1212),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12355_ (.CLK(clknet_leaf_105_clk),
    .D(net2741),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12356_ (.CLK(clknet_leaf_106_clk),
    .D(net2335),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12357_ (.CLK(clknet_leaf_105_clk),
    .D(net2525),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12358_ (.CLK(clknet_leaf_109_clk),
    .D(net774),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12359_ (.CLK(clknet_leaf_111_clk),
    .D(net1217),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12360_ (.CLK(clknet_leaf_109_clk),
    .D(net1107),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12361_ (.CLK(clknet_leaf_109_clk),
    .D(net798),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12362_ (.CLK(clknet_leaf_105_clk),
    .D(net239),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12363_ (.CLK(clknet_leaf_112_clk),
    .D(net1059),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12364_ (.CLK(clknet_leaf_111_clk),
    .D(net1201),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12365_ (.CLK(clknet_leaf_111_clk),
    .D(net466),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12366_ (.CLK(clknet_leaf_74_clk),
    .D(net1147),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12367_ (.CLK(clknet_leaf_74_clk),
    .D(net2827),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12368_ (.CLK(clknet_leaf_74_clk),
    .D(net2762),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12369_ (.CLK(clknet_leaf_115_clk),
    .D(net1359),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12370_ (.CLK(clknet_leaf_115_clk),
    .D(net2943),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12371_ (.CLK(clknet_leaf_115_clk),
    .D(net1394),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12372_ (.CLK(clknet_leaf_115_clk),
    .D(net2849),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12373_ (.CLK(clknet_leaf_115_clk),
    .D(net462),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12374_ (.CLK(clknet_leaf_116_clk),
    .D(net814),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12375_ (.CLK(clknet_leaf_117_clk),
    .D(net2384),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12376_ (.CLK(clknet_leaf_117_clk),
    .D(net1248),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12377_ (.CLK(clknet_leaf_116_clk),
    .D(net1801),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12378_ (.CLK(clknet_leaf_118_clk),
    .D(net438),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _12379_ (.CLK(clknet_leaf_119_clk),
    .D(net503),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _12380_ (.CLK(clknet_leaf_118_clk),
    .D(net2333),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_2 _12381_ (.CLK(clknet_leaf_115_clk),
    .D(_00073_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _12382_ (.CLK(clknet_leaf_116_clk),
    .D(_00074_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12383_ (.CLK(clknet_leaf_116_clk),
    .D(_00075_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12384_ (.CLK(clknet_leaf_111_clk),
    .D(_00076_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12385_ (.CLK(clknet_leaf_116_clk),
    .D(_00077_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12386_ (.CLK(clknet_leaf_116_clk),
    .D(_00078_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12387_ (.CLK(clknet_leaf_116_clk),
    .D(_00079_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12388_ (.CLK(clknet_leaf_115_clk),
    .D(_00080_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ));
 sky130_fd_sc_hd__dfxtp_1 _12389_ (.CLK(clknet_leaf_118_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12390_ (.CLK(clknet_leaf_118_clk),
    .D(net2546),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12391_ (.CLK(clknet_leaf_118_clk),
    .D(net1275),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12392_ (.CLK(clknet_leaf_118_clk),
    .D(net2215),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12393_ (.CLK(clknet_leaf_109_clk),
    .D(_00015_),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _12394_ (.CLK(clknet_leaf_102_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12395_ (.CLK(clknet_leaf_105_clk),
    .D(net2992),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12396_ (.CLK(clknet_leaf_105_clk),
    .D(net3070),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12397_ (.CLK(clknet_leaf_109_clk),
    .D(net3011),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12398_ (.CLK(clknet_leaf_111_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12399_ (.CLK(clknet_leaf_111_clk),
    .D(net3097),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12400_ (.CLK(clknet_leaf_111_clk),
    .D(net3008),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12401_ (.CLK(clknet_leaf_111_clk),
    .D(net3018),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12402_ (.CLK(clknet_leaf_116_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12403_ (.CLK(clknet_leaf_111_clk),
    .D(net2946),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12404_ (.CLK(clknet_leaf_111_clk),
    .D(net3016),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12405_ (.CLK(clknet_leaf_109_clk),
    .D(net2991),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12406_ (.CLK(clknet_leaf_111_clk),
    .D(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12407_ (.CLK(clknet_leaf_111_clk),
    .D(net3129),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12408_ (.CLK(clknet_leaf_108_clk),
    .D(net3126),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12409_ (.CLK(clknet_leaf_108_clk),
    .D(net3127),
    .Q(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12410_ (.CLK(clknet_leaf_130_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12411_ (.CLK(clknet_leaf_130_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12412_ (.CLK(clknet_leaf_108_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12413_ (.CLK(clknet_leaf_109_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12414_ (.CLK(clknet_leaf_132_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12415_ (.CLK(clknet_leaf_107_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12416_ (.CLK(clknet_leaf_132_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12417_ (.CLK(clknet_leaf_132_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12418_ (.CLK(clknet_leaf_129_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12419_ (.CLK(clknet_leaf_130_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12420_ (.CLK(clknet_leaf_130_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12421_ (.CLK(clknet_leaf_129_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12422_ (.CLK(clknet_leaf_131_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12423_ (.CLK(clknet_leaf_132_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12424_ (.CLK(clknet_leaf_132_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12425_ (.CLK(clknet_leaf_133_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12426_ (.CLK(clknet_leaf_128_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12427_ (.CLK(clknet_leaf_130_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12428_ (.CLK(clknet_leaf_130_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12429_ (.CLK(clknet_leaf_130_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12430_ (.CLK(clknet_leaf_133_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12431_ (.CLK(clknet_leaf_133_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12432_ (.CLK(clknet_leaf_133_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12433_ (.CLK(clknet_leaf_133_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12434_ (.CLK(clknet_leaf_128_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12435_ (.CLK(clknet_leaf_128_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12436_ (.CLK(clknet_leaf_128_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12437_ (.CLK(clknet_leaf_128_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12438_ (.CLK(clknet_leaf_133_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12439_ (.CLK(clknet_leaf_134_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12440_ (.CLK(clknet_leaf_134_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12441_ (.CLK(clknet_leaf_134_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12442_ (.CLK(clknet_leaf_123_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12443_ (.CLK(clknet_leaf_123_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12444_ (.CLK(clknet_leaf_122_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12445_ (.CLK(clknet_leaf_124_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12446_ (.CLK(clknet_leaf_123_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12447_ (.CLK(clknet_leaf_123_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12448_ (.CLK(clknet_leaf_123_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12449_ (.CLK(clknet_leaf_123_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12450_ (.CLK(clknet_leaf_124_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12451_ (.CLK(clknet_leaf_129_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12452_ (.CLK(clknet_leaf_128_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12453_ (.CLK(clknet_leaf_124_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12454_ (.CLK(clknet_leaf_119_clk),
    .D(net3272),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12455_ (.CLK(clknet_leaf_119_clk),
    .D(net3235),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12456_ (.CLK(clknet_leaf_117_clk),
    .D(net3254),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12457_ (.CLK(clknet_leaf_130_clk),
    .D(net2450),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12458_ (.CLK(clknet_leaf_131_clk),
    .D(net864),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12459_ (.CLK(clknet_leaf_108_clk),
    .D(net835),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12460_ (.CLK(clknet_leaf_108_clk),
    .D(net530),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12461_ (.CLK(clknet_leaf_132_clk),
    .D(net2357),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12462_ (.CLK(clknet_leaf_132_clk),
    .D(net194),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12463_ (.CLK(clknet_leaf_107_clk),
    .D(net83),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12464_ (.CLK(clknet_leaf_132_clk),
    .D(net1678),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12465_ (.CLK(clknet_leaf_129_clk),
    .D(net974),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12466_ (.CLK(clknet_leaf_130_clk),
    .D(net1472),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12467_ (.CLK(clknet_leaf_130_clk),
    .D(net1648),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12468_ (.CLK(clknet_leaf_110_clk),
    .D(net64),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12469_ (.CLK(clknet_leaf_131_clk),
    .D(net956),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12470_ (.CLK(clknet_leaf_132_clk),
    .D(net2698),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12471_ (.CLK(clknet_leaf_133_clk),
    .D(net489),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12472_ (.CLK(clknet_leaf_133_clk),
    .D(net1172),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12473_ (.CLK(clknet_leaf_131_clk),
    .D(net775),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12474_ (.CLK(clknet_leaf_130_clk),
    .D(net2271),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12475_ (.CLK(clknet_leaf_130_clk),
    .D(net1423),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12476_ (.CLK(clknet_leaf_130_clk),
    .D(net1672),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12477_ (.CLK(clknet_leaf_133_clk),
    .D(net2136),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12478_ (.CLK(clknet_leaf_134_clk),
    .D(net663),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12479_ (.CLK(clknet_leaf_133_clk),
    .D(net2920),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12480_ (.CLK(clknet_leaf_133_clk),
    .D(net1178),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12481_ (.CLK(clknet_leaf_128_clk),
    .D(net2250),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12482_ (.CLK(clknet_leaf_128_clk),
    .D(net1812),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12483_ (.CLK(clknet_leaf_128_clk),
    .D(net976),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12484_ (.CLK(clknet_leaf_128_clk),
    .D(net1020),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12485_ (.CLK(clknet_leaf_135_clk),
    .D(net739),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12486_ (.CLK(clknet_leaf_135_clk),
    .D(net765),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12487_ (.CLK(clknet_leaf_134_clk),
    .D(net1222),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12488_ (.CLK(clknet_leaf_134_clk),
    .D(net1238),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12489_ (.CLK(clknet_leaf_123_clk),
    .D(net2411),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12490_ (.CLK(clknet_leaf_123_clk),
    .D(net1769),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12491_ (.CLK(clknet_leaf_123_clk),
    .D(net265),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12492_ (.CLK(clknet_leaf_124_clk),
    .D(net2674),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12493_ (.CLK(clknet_leaf_123_clk),
    .D(net1722),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12494_ (.CLK(clknet_leaf_117_clk),
    .D(net102),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12495_ (.CLK(clknet_leaf_124_clk),
    .D(net486),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12496_ (.CLK(clknet_leaf_123_clk),
    .D(net1693),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12497_ (.CLK(clknet_leaf_124_clk),
    .D(net1460),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12498_ (.CLK(clknet_leaf_124_clk),
    .D(net84),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12499_ (.CLK(clknet_leaf_128_clk),
    .D(net1595),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12500_ (.CLK(clknet_leaf_124_clk),
    .D(net2412),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12501_ (.CLK(clknet_leaf_117_clk),
    .D(net407),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12502_ (.CLK(clknet_leaf_119_clk),
    .D(net2243),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12503_ (.CLK(clknet_leaf_117_clk),
    .D(net2441),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12504_ (.CLK(clknet_leaf_130_clk),
    .D(net1902),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12505_ (.CLK(clknet_leaf_131_clk),
    .D(net978),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12506_ (.CLK(clknet_leaf_108_clk),
    .D(net834),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12507_ (.CLK(clknet_leaf_108_clk),
    .D(net863),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12508_ (.CLK(clknet_leaf_132_clk),
    .D(net1261),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12509_ (.CLK(clknet_leaf_107_clk),
    .D(net86),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12510_ (.CLK(clknet_leaf_107_clk),
    .D(net1150),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12511_ (.CLK(clknet_leaf_132_clk),
    .D(net1208),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12512_ (.CLK(clknet_leaf_129_clk),
    .D(net836),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12513_ (.CLK(clknet_leaf_130_clk),
    .D(net1292),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12514_ (.CLK(clknet_leaf_130_clk),
    .D(net2257),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12515_ (.CLK(clknet_leaf_129_clk),
    .D(net439),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12516_ (.CLK(clknet_leaf_131_clk),
    .D(net2155),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12517_ (.CLK(clknet_leaf_132_clk),
    .D(net1989),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12518_ (.CLK(clknet_leaf_132_clk),
    .D(net426),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12519_ (.CLK(clknet_leaf_132_clk),
    .D(net409),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12520_ (.CLK(clknet_leaf_131_clk),
    .D(net945),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12521_ (.CLK(clknet_leaf_130_clk),
    .D(net2474),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12522_ (.CLK(clknet_leaf_130_clk),
    .D(net1982),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12523_ (.CLK(clknet_leaf_130_clk),
    .D(net1262),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12524_ (.CLK(clknet_leaf_133_clk),
    .D(net2926),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12525_ (.CLK(clknet_leaf_133_clk),
    .D(net584),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12526_ (.CLK(clknet_leaf_133_clk),
    .D(net2869),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12527_ (.CLK(clknet_leaf_133_clk),
    .D(net2168),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12528_ (.CLK(clknet_leaf_128_clk),
    .D(net1865),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12529_ (.CLK(clknet_leaf_128_clk),
    .D(net964),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12530_ (.CLK(clknet_leaf_128_clk),
    .D(net967),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12531_ (.CLK(clknet_leaf_128_clk),
    .D(net1190),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12532_ (.CLK(clknet_leaf_133_clk),
    .D(net336),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12533_ (.CLK(clknet_leaf_133_clk),
    .D(net358),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12534_ (.CLK(clknet_leaf_134_clk),
    .D(net2513),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12535_ (.CLK(clknet_leaf_134_clk),
    .D(net2626),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12536_ (.CLK(clknet_leaf_123_clk),
    .D(net1652),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12537_ (.CLK(clknet_leaf_123_clk),
    .D(net2809),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12538_ (.CLK(clknet_leaf_122_clk),
    .D(net787),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12539_ (.CLK(clknet_leaf_124_clk),
    .D(net2098),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12540_ (.CLK(clknet_leaf_123_clk),
    .D(net2352),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12541_ (.CLK(clknet_leaf_123_clk),
    .D(net161),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12542_ (.CLK(clknet_leaf_124_clk),
    .D(net2553),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12543_ (.CLK(clknet_leaf_123_clk),
    .D(net1750),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12544_ (.CLK(clknet_leaf_124_clk),
    .D(net2486),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12545_ (.CLK(clknet_leaf_128_clk),
    .D(net238),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12546_ (.CLK(clknet_leaf_128_clk),
    .D(net975),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12547_ (.CLK(clknet_leaf_124_clk),
    .D(net2200),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12548_ (.CLK(clknet_leaf_117_clk),
    .D(net1249),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12549_ (.CLK(clknet_leaf_119_clk),
    .D(net1429),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12550_ (.CLK(clknet_leaf_117_clk),
    .D(net2210),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12551_ (.CLK(clknet_leaf_130_clk),
    .D(net1527),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12552_ (.CLK(clknet_leaf_132_clk),
    .D(net209),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12553_ (.CLK(clknet_leaf_132_clk),
    .D(net152),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12554_ (.CLK(clknet_leaf_132_clk),
    .D(net148),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12555_ (.CLK(clknet_leaf_132_clk),
    .D(net2414),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12556_ (.CLK(clknet_leaf_132_clk),
    .D(net215),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12557_ (.CLK(clknet_leaf_132_clk),
    .D(net217),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12558_ (.CLK(clknet_leaf_132_clk),
    .D(net1904),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12559_ (.CLK(clknet_leaf_129_clk),
    .D(net1070),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12560_ (.CLK(clknet_leaf_130_clk),
    .D(net1311),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12561_ (.CLK(clknet_leaf_130_clk),
    .D(net1609),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12562_ (.CLK(clknet_leaf_129_clk),
    .D(net825),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12563_ (.CLK(clknet_leaf_132_clk),
    .D(net195),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12564_ (.CLK(clknet_leaf_132_clk),
    .D(net2531),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12565_ (.CLK(clknet_leaf_132_clk),
    .D(net2005),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12566_ (.CLK(clknet_leaf_133_clk),
    .D(net699),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _12567_ (.CLK(clknet_leaf_131_clk),
    .D(net857),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12568_ (.CLK(clknet_leaf_130_clk),
    .D(net2223),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12569_ (.CLK(clknet_leaf_130_clk),
    .D(net1232),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12570_ (.CLK(clknet_leaf_130_clk),
    .D(net2278),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _12571_ (.CLK(clknet_leaf_133_clk),
    .D(net2848),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12572_ (.CLK(clknet_leaf_133_clk),
    .D(net2944),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12573_ (.CLK(clknet_leaf_133_clk),
    .D(net2942),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12574_ (.CLK(clknet_leaf_133_clk),
    .D(net2400),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12575_ (.CLK(clknet_leaf_128_clk),
    .D(net1026),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12576_ (.CLK(clknet_leaf_131_clk),
    .D(net786),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12577_ (.CLK(clknet_leaf_131_clk),
    .D(net785),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12578_ (.CLK(clknet_leaf_128_clk),
    .D(net2011),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12579_ (.CLK(clknet_leaf_133_clk),
    .D(net2493),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_2 _12580_ (.CLK(clknet_leaf_133_clk),
    .D(net1220),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12581_ (.CLK(clknet_leaf_134_clk),
    .D(net1252),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12582_ (.CLK(clknet_leaf_134_clk),
    .D(net2551),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12583_ (.CLK(clknet_leaf_123_clk),
    .D(net1299),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12584_ (.CLK(clknet_leaf_129_clk),
    .D(net700),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12585_ (.CLK(clknet_leaf_123_clk),
    .D(net275),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12586_ (.CLK(clknet_leaf_124_clk),
    .D(net2590),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12587_ (.CLK(clknet_leaf_123_clk),
    .D(net1732),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12588_ (.CLK(clknet_leaf_123_clk),
    .D(net1860),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12589_ (.CLK(clknet_leaf_124_clk),
    .D(net2902),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12590_ (.CLK(clknet_leaf_124_clk),
    .D(net474),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12591_ (.CLK(clknet_leaf_124_clk),
    .D(net2932),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12592_ (.CLK(clknet_leaf_129_clk),
    .D(net1863),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12593_ (.CLK(clknet_leaf_128_clk),
    .D(net1805),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12594_ (.CLK(clknet_leaf_124_clk),
    .D(net1518),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12595_ (.CLK(clknet_leaf_117_clk),
    .D(net2381),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _12596_ (.CLK(clknet_leaf_119_clk),
    .D(net1187),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _12597_ (.CLK(clknet_leaf_117_clk),
    .D(net1853),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _12598_ (.CLK(clknet_leaf_129_clk),
    .D(_00081_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _12599_ (.CLK(clknet_leaf_124_clk),
    .D(_00082_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12600_ (.CLK(clknet_leaf_123_clk),
    .D(_00083_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12601_ (.CLK(clknet_leaf_123_clk),
    .D(_00084_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12602_ (.CLK(clknet_leaf_129_clk),
    .D(_00085_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12603_ (.CLK(clknet_leaf_129_clk),
    .D(_00086_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12604_ (.CLK(clknet_leaf_129_clk),
    .D(_00087_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _12605_ (.CLK(clknet_leaf_168_clk),
    .D(_00088_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ));
 sky130_fd_sc_hd__dfxtp_1 _12606_ (.CLK(clknet_leaf_117_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12607_ (.CLK(clknet_leaf_117_clk),
    .D(net1993),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12608_ (.CLK(clknet_leaf_117_clk),
    .D(net2399),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12609_ (.CLK(clknet_leaf_117_clk),
    .D(net2386),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12610_ (.CLK(clknet_leaf_134_clk),
    .D(_00008_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _12611_ (.CLK(clknet_leaf_124_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12612_ (.CLK(clknet_leaf_134_clk),
    .D(net3080),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12613_ (.CLK(clknet_leaf_131_clk),
    .D(net3099),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12614_ (.CLK(clknet_leaf_131_clk),
    .D(net3032),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12615_ (.CLK(clknet_leaf_124_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12616_ (.CLK(clknet_leaf_132_clk),
    .D(net3075),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12617_ (.CLK(clknet_leaf_131_clk),
    .D(net3096),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12618_ (.CLK(clknet_leaf_131_clk),
    .D(net3056),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12619_ (.CLK(clknet_leaf_124_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12620_ (.CLK(clknet_leaf_131_clk),
    .D(net3110),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12621_ (.CLK(clknet_leaf_134_clk),
    .D(net2948),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12622_ (.CLK(clknet_leaf_134_clk),
    .D(net3066),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12623_ (.CLK(clknet_leaf_128_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12624_ (.CLK(clknet_leaf_131_clk),
    .D(net3135),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12625_ (.CLK(clknet_leaf_134_clk),
    .D(net2977),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12626_ (.CLK(clknet_leaf_133_clk),
    .D(net3036),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12627_ (.CLK(clknet_leaf_134_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12628_ (.CLK(clknet_leaf_135_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12629_ (.CLK(clknet_leaf_135_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12630_ (.CLK(clknet_leaf_135_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12631_ (.CLK(clknet_leaf_136_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12632_ (.CLK(clknet_leaf_142_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12633_ (.CLK(clknet_leaf_136_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12634_ (.CLK(clknet_leaf_142_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12635_ (.CLK(clknet_leaf_127_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12636_ (.CLK(clknet_leaf_127_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12637_ (.CLK(clknet_leaf_137_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12638_ (.CLK(clknet_leaf_127_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12639_ (.CLK(clknet_leaf_135_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12640_ (.CLK(clknet_leaf_135_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12641_ (.CLK(clknet_leaf_134_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12642_ (.CLK(clknet_leaf_136_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12643_ (.CLK(clknet_leaf_128_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12644_ (.CLK(clknet_leaf_138_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12645_ (.CLK(clknet_leaf_126_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12646_ (.CLK(clknet_leaf_127_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12647_ (.CLK(clknet_leaf_136_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12648_ (.CLK(clknet_leaf_136_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12649_ (.CLK(clknet_leaf_137_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12650_ (.CLK(clknet_leaf_137_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12651_ (.CLK(clknet_leaf_138_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12652_ (.CLK(clknet_leaf_139_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12653_ (.CLK(clknet_leaf_139_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12654_ (.CLK(clknet_leaf_138_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12655_ (.CLK(clknet_leaf_141_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12656_ (.CLK(clknet_leaf_141_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12657_ (.CLK(clknet_leaf_140_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12658_ (.CLK(clknet_leaf_141_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12659_ (.CLK(clknet_leaf_125_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12660_ (.CLK(clknet_leaf_125_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12661_ (.CLK(clknet_leaf_125_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12662_ (.CLK(clknet_leaf_125_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12663_ (.CLK(clknet_leaf_125_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12664_ (.CLK(clknet_leaf_162_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12665_ (.CLK(clknet_leaf_126_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12666_ (.CLK(clknet_leaf_126_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12667_ (.CLK(clknet_leaf_126_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12668_ (.CLK(clknet_leaf_126_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12669_ (.CLK(clknet_leaf_138_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12670_ (.CLK(clknet_leaf_126_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12671_ (.CLK(clknet_leaf_119_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12672_ (.CLK(clknet_leaf_119_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12673_ (.CLK(clknet_leaf_119_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12674_ (.CLK(clknet_leaf_134_clk),
    .D(net2460),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12675_ (.CLK(clknet_leaf_135_clk),
    .D(net1395),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12676_ (.CLK(clknet_leaf_134_clk),
    .D(net323),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12677_ (.CLK(clknet_leaf_135_clk),
    .D(net2358),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12678_ (.CLK(clknet_leaf_136_clk),
    .D(net1586),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12679_ (.CLK(clknet_leaf_142_clk),
    .D(net1231),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12680_ (.CLK(clknet_leaf_136_clk),
    .D(net1017),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12681_ (.CLK(clknet_leaf_142_clk),
    .D(net2405),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12682_ (.CLK(clknet_leaf_127_clk),
    .D(net869),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12683_ (.CLK(clknet_leaf_127_clk),
    .D(net860),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12684_ (.CLK(clknet_leaf_137_clk),
    .D(net2368),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12685_ (.CLK(clknet_leaf_127_clk),
    .D(net902),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12686_ (.CLK(clknet_leaf_135_clk),
    .D(net1164),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12687_ (.CLK(clknet_leaf_135_clk),
    .D(net1811),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12688_ (.CLK(clknet_leaf_137_clk),
    .D(net533),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12689_ (.CLK(clknet_leaf_136_clk),
    .D(net2236),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12690_ (.CLK(clknet_leaf_127_clk),
    .D(net762),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12691_ (.CLK(clknet_leaf_138_clk),
    .D(net999),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12692_ (.CLK(clknet_leaf_137_clk),
    .D(net633),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12693_ (.CLK(clknet_leaf_137_clk),
    .D(net225),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12694_ (.CLK(clknet_leaf_136_clk),
    .D(net1029),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12695_ (.CLK(clknet_leaf_136_clk),
    .D(net1772),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12696_ (.CLK(clknet_leaf_137_clk),
    .D(net2121),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12697_ (.CLK(clknet_leaf_134_clk),
    .D(net655),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12698_ (.CLK(clknet_leaf_138_clk),
    .D(net2319),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12699_ (.CLK(clknet_leaf_139_clk),
    .D(net2635),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12700_ (.CLK(clknet_leaf_139_clk),
    .D(net1230),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12701_ (.CLK(clknet_leaf_138_clk),
    .D(net1176),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12702_ (.CLK(clknet_leaf_141_clk),
    .D(net1475),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12703_ (.CLK(clknet_leaf_141_clk),
    .D(net1325),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12704_ (.CLK(clknet_leaf_141_clk),
    .D(net604),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12705_ (.CLK(clknet_leaf_141_clk),
    .D(net1762),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12706_ (.CLK(clknet_leaf_124_clk),
    .D(net297),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12707_ (.CLK(clknet_leaf_125_clk),
    .D(net2102),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12708_ (.CLK(clknet_leaf_124_clk),
    .D(net319),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12709_ (.CLK(clknet_leaf_125_clk),
    .D(net2208),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12710_ (.CLK(clknet_leaf_162_clk),
    .D(net473),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12711_ (.CLK(clknet_leaf_162_clk),
    .D(net2578),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12712_ (.CLK(clknet_leaf_126_clk),
    .D(net2833),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12713_ (.CLK(clknet_leaf_126_clk),
    .D(net1833),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12714_ (.CLK(clknet_leaf_126_clk),
    .D(net2691),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12715_ (.CLK(clknet_leaf_126_clk),
    .D(net2494),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12716_ (.CLK(clknet_leaf_138_clk),
    .D(net2797),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12717_ (.CLK(clknet_leaf_126_clk),
    .D(net1976),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12718_ (.CLK(clknet_leaf_120_clk),
    .D(net160),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12719_ (.CLK(clknet_leaf_120_clk),
    .D(net156),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12720_ (.CLK(clknet_leaf_117_clk),
    .D(net339),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12721_ (.CLK(clknet_leaf_134_clk),
    .D(net1565),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12722_ (.CLK(clknet_leaf_135_clk),
    .D(net1963),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12723_ (.CLK(clknet_leaf_135_clk),
    .D(net679),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12724_ (.CLK(clknet_leaf_135_clk),
    .D(net1910),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12725_ (.CLK(clknet_leaf_136_clk),
    .D(net2672),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12726_ (.CLK(clknet_leaf_136_clk),
    .D(net747),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12727_ (.CLK(clknet_leaf_136_clk),
    .D(net1857),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12728_ (.CLK(clknet_leaf_142_clk),
    .D(net2314),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12729_ (.CLK(clknet_leaf_137_clk),
    .D(net242),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12730_ (.CLK(clknet_leaf_127_clk),
    .D(net2330),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12731_ (.CLK(clknet_leaf_137_clk),
    .D(net1483),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12732_ (.CLK(clknet_leaf_137_clk),
    .D(net229),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12733_ (.CLK(clknet_leaf_135_clk),
    .D(net2186),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12734_ (.CLK(clknet_leaf_135_clk),
    .D(net1946),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12735_ (.CLK(clknet_leaf_134_clk),
    .D(net596),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12736_ (.CLK(clknet_leaf_135_clk),
    .D(net271),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12737_ (.CLK(clknet_leaf_127_clk),
    .D(net851),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12738_ (.CLK(clknet_leaf_138_clk),
    .D(net1303),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12739_ (.CLK(clknet_leaf_137_clk),
    .D(net2069),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12740_ (.CLK(clknet_leaf_137_clk),
    .D(net2699),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12741_ (.CLK(clknet_leaf_136_clk),
    .D(net2088),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12742_ (.CLK(clknet_leaf_136_clk),
    .D(net1753),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12743_ (.CLK(clknet_leaf_137_clk),
    .D(net2756),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12744_ (.CLK(clknet_leaf_137_clk),
    .D(net465),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12745_ (.CLK(clknet_leaf_138_clk),
    .D(net2515),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12746_ (.CLK(clknet_leaf_139_clk),
    .D(net2063),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12747_ (.CLK(clknet_leaf_139_clk),
    .D(net2713),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12748_ (.CLK(clknet_leaf_138_clk),
    .D(net1093),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12749_ (.CLK(clknet_leaf_141_clk),
    .D(net1838),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12750_ (.CLK(clknet_leaf_141_clk),
    .D(net2489),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12751_ (.CLK(clknet_leaf_141_clk),
    .D(net1647),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12752_ (.CLK(clknet_leaf_141_clk),
    .D(net2225),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12753_ (.CLK(clknet_leaf_124_clk),
    .D(net2638),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12754_ (.CLK(clknet_leaf_125_clk),
    .D(net1675),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12755_ (.CLK(clknet_leaf_125_clk),
    .D(net703),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12756_ (.CLK(clknet_leaf_125_clk),
    .D(net1080),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12757_ (.CLK(clknet_leaf_125_clk),
    .D(net569),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12758_ (.CLK(clknet_leaf_162_clk),
    .D(net1388),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12759_ (.CLK(clknet_leaf_126_clk),
    .D(net2140),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12760_ (.CLK(clknet_leaf_125_clk),
    .D(net145),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12761_ (.CLK(clknet_leaf_126_clk),
    .D(net2117),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12762_ (.CLK(clknet_leaf_126_clk),
    .D(net2851),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12763_ (.CLK(clknet_leaf_138_clk),
    .D(net2722),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12764_ (.CLK(clknet_leaf_126_clk),
    .D(net2449),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12765_ (.CLK(clknet_leaf_119_clk),
    .D(net110),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12766_ (.CLK(clknet_leaf_119_clk),
    .D(net105),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12767_ (.CLK(clknet_leaf_122_clk),
    .D(net172),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12768_ (.CLK(clknet_leaf_134_clk),
    .D(net2402),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12769_ (.CLK(clknet_leaf_135_clk),
    .D(net1337),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12770_ (.CLK(clknet_leaf_135_clk),
    .D(net1437),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12771_ (.CLK(clknet_leaf_135_clk),
    .D(net1978),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12772_ (.CLK(clknet_leaf_136_clk),
    .D(net2879),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12773_ (.CLK(clknet_leaf_142_clk),
    .D(net631),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12774_ (.CLK(clknet_leaf_136_clk),
    .D(net1570),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12775_ (.CLK(clknet_leaf_142_clk),
    .D(net2884),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12776_ (.CLK(clknet_leaf_137_clk),
    .D(net2111),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12777_ (.CLK(clknet_leaf_127_clk),
    .D(net1060),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12778_ (.CLK(clknet_leaf_137_clk),
    .D(net2658),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12779_ (.CLK(clknet_leaf_137_clk),
    .D(net2908),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12780_ (.CLK(clknet_leaf_135_clk),
    .D(net1841),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12781_ (.CLK(clknet_leaf_136_clk),
    .D(net154),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12782_ (.CLK(clknet_leaf_134_clk),
    .D(net2079),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12783_ (.CLK(clknet_leaf_135_clk),
    .D(net2146),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _12784_ (.CLK(clknet_leaf_127_clk),
    .D(net884),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12785_ (.CLK(clknet_leaf_137_clk),
    .D(net212),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12786_ (.CLK(clknet_leaf_138_clk),
    .D(net164),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12787_ (.CLK(clknet_leaf_137_clk),
    .D(net1977),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _12788_ (.CLK(clknet_leaf_136_clk),
    .D(net2585),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12789_ (.CLK(clknet_leaf_136_clk),
    .D(net2040),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12790_ (.CLK(clknet_leaf_137_clk),
    .D(net1640),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12791_ (.CLK(clknet_leaf_134_clk),
    .D(net672),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12792_ (.CLK(clknet_leaf_138_clk),
    .D(net1276),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12793_ (.CLK(clknet_leaf_139_clk),
    .D(net1120),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12794_ (.CLK(clknet_leaf_139_clk),
    .D(net2706),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12795_ (.CLK(clknet_leaf_138_clk),
    .D(net981),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12796_ (.CLK(clknet_leaf_142_clk),
    .D(net435),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12797_ (.CLK(clknet_leaf_142_clk),
    .D(net757),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12798_ (.CLK(clknet_leaf_141_clk),
    .D(net2700),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12799_ (.CLK(clknet_leaf_141_clk),
    .D(net2538),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12800_ (.CLK(clknet_leaf_125_clk),
    .D(net806),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12801_ (.CLK(clknet_leaf_125_clk),
    .D(net2109),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12802_ (.CLK(clknet_leaf_124_clk),
    .D(net308),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12803_ (.CLK(clknet_leaf_125_clk),
    .D(net2313),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12804_ (.CLK(clknet_leaf_125_clk),
    .D(net2191),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12805_ (.CLK(clknet_leaf_125_clk),
    .D(net499),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12806_ (.CLK(clknet_leaf_126_clk),
    .D(net2858),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12807_ (.CLK(clknet_leaf_126_clk),
    .D(net181),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12808_ (.CLK(clknet_leaf_138_clk),
    .D(net168),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12809_ (.CLK(clknet_leaf_126_clk),
    .D(net2832),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12810_ (.CLK(clknet_leaf_138_clk),
    .D(net1061),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12811_ (.CLK(clknet_leaf_138_clk),
    .D(net187),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12812_ (.CLK(clknet_leaf_121_clk),
    .D(net159),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _12813_ (.CLK(clknet_leaf_119_clk),
    .D(net2075),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _12814_ (.CLK(clknet_leaf_117_clk),
    .D(net90),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _12815_ (.CLK(clknet_leaf_127_clk),
    .D(_00089_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _12816_ (.CLK(clknet_leaf_127_clk),
    .D(_00090_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12817_ (.CLK(clknet_leaf_127_clk),
    .D(_00091_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12818_ (.CLK(clknet_leaf_127_clk),
    .D(_00092_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12819_ (.CLK(clknet_leaf_126_clk),
    .D(_00093_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12820_ (.CLK(clknet_leaf_127_clk),
    .D(_00094_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12821_ (.CLK(clknet_leaf_127_clk),
    .D(_00095_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12822_ (.CLK(clknet_leaf_122_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12823_ (.CLK(clknet_leaf_122_clk),
    .D(net1119),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12824_ (.CLK(clknet_leaf_122_clk),
    .D(net1735),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12825_ (.CLK(clknet_leaf_123_clk),
    .D(net291),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12826_ (.CLK(clknet_leaf_137_clk),
    .D(_00009_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _12827_ (.CLK(clknet_leaf_125_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12828_ (.CLK(clknet_leaf_136_clk),
    .D(net2995),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12829_ (.CLK(clknet_leaf_137_clk),
    .D(net2957),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12830_ (.CLK(clknet_leaf_137_clk),
    .D(net3052),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12831_ (.CLK(clknet_leaf_126_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12832_ (.CLK(clknet_leaf_138_clk),
    .D(net3014),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12833_ (.CLK(clknet_leaf_141_clk),
    .D(net2985),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12834_ (.CLK(clknet_leaf_139_clk),
    .D(net2999),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12835_ (.CLK(clknet_leaf_126_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12836_ (.CLK(clknet_leaf_138_clk),
    .D(net2996),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12837_ (.CLK(clknet_leaf_138_clk),
    .D(net3109),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12838_ (.CLK(clknet_leaf_138_clk),
    .D(net3112),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12839_ (.CLK(clknet_leaf_126_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12840_ (.CLK(clknet_leaf_136_clk),
    .D(net2997),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12841_ (.CLK(clknet_leaf_136_clk),
    .D(net3122),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12842_ (.CLK(clknet_leaf_137_clk),
    .D(net2969),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12843_ (.CLK(clknet_leaf_142_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12844_ (.CLK(clknet_leaf_142_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12845_ (.CLK(clknet_leaf_141_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12846_ (.CLK(clknet_leaf_141_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12847_ (.CLK(clknet_leaf_142_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12848_ (.CLK(clknet_leaf_143_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12849_ (.CLK(clknet_leaf_143_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12850_ (.CLK(clknet_leaf_143_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12851_ (.CLK(clknet_leaf_139_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12852_ (.CLK(clknet_leaf_139_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12853_ (.CLK(clknet_leaf_139_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12854_ (.CLK(clknet_leaf_140_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12855_ (.CLK(clknet_leaf_141_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12856_ (.CLK(clknet_leaf_141_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12857_ (.CLK(clknet_leaf_140_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12858_ (.CLK(clknet_leaf_140_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12859_ (.CLK(clknet_leaf_146_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12860_ (.CLK(clknet_leaf_148_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12861_ (.CLK(clknet_leaf_147_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12862_ (.CLK(clknet_leaf_148_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12863_ (.CLK(clknet_leaf_144_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12864_ (.CLK(clknet_leaf_144_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12865_ (.CLK(clknet_leaf_144_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12866_ (.CLK(clknet_leaf_144_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12867_ (.CLK(clknet_leaf_147_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12868_ (.CLK(clknet_leaf_147_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12869_ (.CLK(clknet_leaf_147_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12870_ (.CLK(clknet_leaf_148_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12871_ (.CLK(clknet_leaf_145_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12872_ (.CLK(clknet_leaf_145_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12873_ (.CLK(clknet_leaf_145_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12874_ (.CLK(clknet_leaf_147_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12875_ (.CLK(clknet_leaf_161_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12876_ (.CLK(clknet_leaf_161_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12877_ (.CLK(clknet_leaf_161_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12878_ (.CLK(clknet_leaf_161_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12879_ (.CLK(clknet_leaf_161_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12880_ (.CLK(clknet_leaf_149_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12881_ (.CLK(clknet_leaf_161_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12882_ (.CLK(clknet_leaf_139_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12883_ (.CLK(clknet_leaf_139_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12884_ (.CLK(clknet_leaf_149_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12885_ (.CLK(clknet_leaf_149_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12886_ (.CLK(clknet_leaf_149_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12887_ (.CLK(clknet_leaf_121_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12888_ (.CLK(clknet_leaf_120_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12889_ (.CLK(clknet_leaf_122_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12890_ (.CLK(clknet_leaf_142_clk),
    .D(net2719),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12891_ (.CLK(clknet_leaf_142_clk),
    .D(net1194),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12892_ (.CLK(clknet_leaf_141_clk),
    .D(net1228),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12893_ (.CLK(clknet_leaf_142_clk),
    .D(net634),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12894_ (.CLK(clknet_leaf_142_clk),
    .D(net1714),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12895_ (.CLK(clknet_leaf_143_clk),
    .D(net993),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12896_ (.CLK(clknet_leaf_143_clk),
    .D(net2526),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12897_ (.CLK(clknet_leaf_143_clk),
    .D(net1013),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12898_ (.CLK(clknet_leaf_140_clk),
    .D(net416),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12899_ (.CLK(clknet_leaf_139_clk),
    .D(net2630),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12900_ (.CLK(clknet_leaf_140_clk),
    .D(net391),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12901_ (.CLK(clknet_leaf_140_clk),
    .D(net1361),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12902_ (.CLK(clknet_leaf_141_clk),
    .D(net1258),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12903_ (.CLK(clknet_leaf_141_clk),
    .D(net1888),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12904_ (.CLK(clknet_leaf_143_clk),
    .D(net620),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12905_ (.CLK(clknet_leaf_143_clk),
    .D(net713),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12906_ (.CLK(clknet_leaf_146_clk),
    .D(net1592),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12907_ (.CLK(clknet_leaf_147_clk),
    .D(net201),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12908_ (.CLK(clknet_leaf_147_clk),
    .D(net2852),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12909_ (.CLK(clknet_leaf_140_clk),
    .D(net192),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12910_ (.CLK(clknet_leaf_144_clk),
    .D(net957),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12911_ (.CLK(clknet_leaf_144_clk),
    .D(net2826),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12912_ (.CLK(clknet_leaf_144_clk),
    .D(net1459),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12913_ (.CLK(clknet_leaf_143_clk),
    .D(net276),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12914_ (.CLK(clknet_leaf_148_clk),
    .D(net969),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12915_ (.CLK(clknet_leaf_147_clk),
    .D(net1618),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12916_ (.CLK(clknet_leaf_147_clk),
    .D(net2940),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12917_ (.CLK(clknet_leaf_140_clk),
    .D(net200),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12918_ (.CLK(clknet_leaf_145_clk),
    .D(net840),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12919_ (.CLK(clknet_leaf_145_clk),
    .D(net901),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12920_ (.CLK(clknet_leaf_145_clk),
    .D(net1016),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12921_ (.CLK(clknet_leaf_145_clk),
    .D(net1087),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12922_ (.CLK(clknet_leaf_161_clk),
    .D(net1957),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12923_ (.CLK(clknet_leaf_126_clk),
    .D(net370),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12924_ (.CLK(clknet_leaf_161_clk),
    .D(net1630),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12925_ (.CLK(clknet_leaf_161_clk),
    .D(net1992),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12926_ (.CLK(clknet_leaf_161_clk),
    .D(net2841),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12927_ (.CLK(clknet_leaf_139_clk),
    .D(net218),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12928_ (.CLK(clknet_leaf_149_clk),
    .D(net537),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12929_ (.CLK(clknet_leaf_139_clk),
    .D(net1551),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12930_ (.CLK(clknet_leaf_139_clk),
    .D(net1790),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12931_ (.CLK(clknet_leaf_149_clk),
    .D(net2746),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12932_ (.CLK(clknet_leaf_149_clk),
    .D(net2503),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12933_ (.CLK(clknet_leaf_149_clk),
    .D(net2561),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12934_ (.CLK(clknet_leaf_121_clk),
    .D(net2656),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12935_ (.CLK(clknet_leaf_120_clk),
    .D(net1366),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12936_ (.CLK(clknet_leaf_122_clk),
    .D(net1757),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12937_ (.CLK(clknet_leaf_142_clk),
    .D(net2938),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12938_ (.CLK(clknet_leaf_142_clk),
    .D(net1350),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12939_ (.CLK(clknet_leaf_142_clk),
    .D(net463),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12940_ (.CLK(clknet_leaf_142_clk),
    .D(net2856),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12941_ (.CLK(clknet_leaf_143_clk),
    .D(net691),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12942_ (.CLK(clknet_leaf_143_clk),
    .D(net2748),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12943_ (.CLK(clknet_leaf_143_clk),
    .D(net2702),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12944_ (.CLK(clknet_leaf_143_clk),
    .D(net1851),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12945_ (.CLK(clknet_leaf_140_clk),
    .D(net2776),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12946_ (.CLK(clknet_leaf_140_clk),
    .D(net419),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12947_ (.CLK(clknet_leaf_140_clk),
    .D(net1918),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12948_ (.CLK(clknet_leaf_140_clk),
    .D(net1661),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12949_ (.CLK(clknet_leaf_141_clk),
    .D(net2066),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12950_ (.CLK(clknet_leaf_141_clk),
    .D(net1850),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12951_ (.CLK(clknet_leaf_143_clk),
    .D(net1843),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12952_ (.CLK(clknet_leaf_140_clk),
    .D(net334),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12953_ (.CLK(clknet_leaf_146_clk),
    .D(net1547),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _12954_ (.CLK(clknet_leaf_147_clk),
    .D(net1322),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _12955_ (.CLK(clknet_leaf_147_clk),
    .D(net1728),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _12956_ (.CLK(clknet_leaf_140_clk),
    .D(net1364),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _12957_ (.CLK(clknet_leaf_144_clk),
    .D(net950),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _12958_ (.CLK(clknet_leaf_144_clk),
    .D(net2422),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _12959_ (.CLK(clknet_leaf_144_clk),
    .D(net1260),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _12960_ (.CLK(clknet_leaf_144_clk),
    .D(net753),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _12961_ (.CLK(clknet_leaf_147_clk),
    .D(net203),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _12962_ (.CLK(clknet_leaf_147_clk),
    .D(net1464),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _12963_ (.CLK(clknet_leaf_147_clk),
    .D(net2356),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _12964_ (.CLK(clknet_leaf_140_clk),
    .D(net2825),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _12965_ (.CLK(clknet_leaf_145_clk),
    .D(net2130),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _12966_ (.CLK(clknet_leaf_145_clk),
    .D(net2221),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _12967_ (.CLK(clknet_leaf_145_clk),
    .D(net2184),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _12968_ (.CLK(clknet_leaf_145_clk),
    .D(net852),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _12969_ (.CLK(clknet_leaf_161_clk),
    .D(net2428),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _12970_ (.CLK(clknet_leaf_161_clk),
    .D(net96),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _12971_ (.CLK(clknet_leaf_161_clk),
    .D(net1526),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _12972_ (.CLK(clknet_leaf_161_clk),
    .D(net2897),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _12973_ (.CLK(clknet_leaf_161_clk),
    .D(net1512),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _12974_ (.CLK(clknet_leaf_139_clk),
    .D(net1911),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _12975_ (.CLK(clknet_leaf_149_clk),
    .D(net2559),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _12976_ (.CLK(clknet_leaf_139_clk),
    .D(net1737),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _12977_ (.CLK(clknet_leaf_139_clk),
    .D(net1173),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _12978_ (.CLK(clknet_leaf_149_clk),
    .D(net2274),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _12979_ (.CLK(clknet_leaf_149_clk),
    .D(net2249),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _12980_ (.CLK(clknet_leaf_149_clk),
    .D(net2752),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _12981_ (.CLK(clknet_leaf_121_clk),
    .D(net1265),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _12982_ (.CLK(clknet_leaf_120_clk),
    .D(net1374),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _12983_ (.CLK(clknet_leaf_122_clk),
    .D(net1167),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _12984_ (.CLK(clknet_leaf_142_clk),
    .D(net2880),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12985_ (.CLK(clknet_leaf_142_clk),
    .D(net2459),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12986_ (.CLK(clknet_leaf_141_clk),
    .D(net602),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12987_ (.CLK(clknet_leaf_142_clk),
    .D(net2881),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12988_ (.CLK(clknet_leaf_143_clk),
    .D(net2549),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12989_ (.CLK(clknet_leaf_143_clk),
    .D(net2562),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12990_ (.CLK(clknet_leaf_143_clk),
    .D(net2306),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12991_ (.CLK(clknet_leaf_143_clk),
    .D(net2031),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12992_ (.CLK(clknet_leaf_140_clk),
    .D(net2657),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12993_ (.CLK(clknet_leaf_140_clk),
    .D(net1357),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12994_ (.CLK(clknet_leaf_140_clk),
    .D(net1379),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12995_ (.CLK(clknet_leaf_140_clk),
    .D(net1398),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12996_ (.CLK(clknet_leaf_141_clk),
    .D(net2500),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12997_ (.CLK(clknet_leaf_142_clk),
    .D(net498),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12998_ (.CLK(clknet_leaf_142_clk),
    .D(net355),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12999_ (.CLK(clknet_leaf_143_clk),
    .D(net618),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13000_ (.CLK(clknet_leaf_146_clk),
    .D(net1030),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13001_ (.CLK(clknet_leaf_147_clk),
    .D(net1244),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13002_ (.CLK(clknet_leaf_147_clk),
    .D(net2846),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13003_ (.CLK(clknet_leaf_140_clk),
    .D(net1681),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13004_ (.CLK(clknet_leaf_144_clk),
    .D(net916),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13005_ (.CLK(clknet_leaf_144_clk),
    .D(net1301),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13006_ (.CLK(clknet_leaf_143_clk),
    .D(net299),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13007_ (.CLK(clknet_leaf_144_clk),
    .D(net1372),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13008_ (.CLK(clknet_leaf_140_clk),
    .D(net411),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13009_ (.CLK(clknet_leaf_147_clk),
    .D(net1264),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13010_ (.CLK(clknet_leaf_147_clk),
    .D(net2936),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13011_ (.CLK(clknet_leaf_140_clk),
    .D(net1369),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13012_ (.CLK(clknet_leaf_144_clk),
    .D(net279),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13013_ (.CLK(clknet_leaf_145_clk),
    .D(net839),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13014_ (.CLK(clknet_leaf_145_clk),
    .D(net848),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13015_ (.CLK(clknet_leaf_145_clk),
    .D(net2738),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13016_ (.CLK(clknet_leaf_161_clk),
    .D(net1698),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13017_ (.CLK(clknet_leaf_126_clk),
    .D(net368),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13018_ (.CLK(clknet_leaf_161_clk),
    .D(net1699),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13019_ (.CLK(clknet_leaf_161_clk),
    .D(net2255),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13020_ (.CLK(clknet_leaf_149_clk),
    .D(net719),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13021_ (.CLK(clknet_leaf_139_clk),
    .D(net1953),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13022_ (.CLK(clknet_leaf_139_clk),
    .D(net224),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13023_ (.CLK(clknet_leaf_139_clk),
    .D(net2913),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13024_ (.CLK(clknet_leaf_139_clk),
    .D(net2263),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13025_ (.CLK(clknet_leaf_149_clk),
    .D(net1799),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13026_ (.CLK(clknet_leaf_149_clk),
    .D(net2560),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13027_ (.CLK(clknet_leaf_149_clk),
    .D(net2268),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13028_ (.CLK(clknet_leaf_121_clk),
    .D(net1725),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _13029_ (.CLK(clknet_leaf_121_clk),
    .D(net585),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _13030_ (.CLK(clknet_leaf_123_clk),
    .D(net286),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _13031_ (.CLK(clknet_leaf_149_clk),
    .D(_00096_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _13032_ (.CLK(clknet_leaf_149_clk),
    .D(net3209),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13033_ (.CLK(clknet_leaf_148_clk),
    .D(_00098_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13034_ (.CLK(clknet_leaf_148_clk),
    .D(_00099_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13035_ (.CLK(clknet_leaf_148_clk),
    .D(_00100_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13036_ (.CLK(clknet_leaf_148_clk),
    .D(_00101_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13037_ (.CLK(clknet_leaf_148_clk),
    .D(_00102_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13038_ (.CLK(clknet_leaf_122_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13039_ (.CLK(clknet_leaf_122_clk),
    .D(net1126),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13040_ (.CLK(clknet_leaf_122_clk),
    .D(net2628),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13041_ (.CLK(clknet_leaf_123_clk),
    .D(net353),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13042_ (.CLK(clknet_leaf_140_clk),
    .D(_00010_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _13043_ (.CLK(clknet_leaf_126_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13044_ (.CLK(clknet_leaf_144_clk),
    .D(net3119),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13045_ (.CLK(clknet_leaf_145_clk),
    .D(net3005),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13046_ (.CLK(clknet_leaf_145_clk),
    .D(net3084),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13047_ (.CLK(clknet_leaf_148_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13048_ (.CLK(clknet_leaf_144_clk),
    .D(net3072),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13049_ (.CLK(clknet_leaf_144_clk),
    .D(net3076),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13050_ (.CLK(clknet_leaf_144_clk),
    .D(net3054),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13051_ (.CLK(clknet_leaf_148_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13052_ (.CLK(clknet_leaf_147_clk),
    .D(net2980),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13053_ (.CLK(clknet_leaf_147_clk),
    .D(net3046),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13054_ (.CLK(clknet_leaf_140_clk),
    .D(net2974),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13055_ (.CLK(clknet_leaf_149_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13056_ (.CLK(clknet_leaf_143_clk),
    .D(net3081),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13057_ (.CLK(clknet_leaf_143_clk),
    .D(net3120),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13058_ (.CLK(clknet_leaf_143_clk),
    .D(net3118),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13059_ (.CLK(clknet_leaf_152_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13060_ (.CLK(clknet_leaf_153_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13061_ (.CLK(clknet_leaf_153_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13062_ (.CLK(clknet_leaf_153_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13063_ (.CLK(clknet_leaf_152_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13064_ (.CLK(clknet_leaf_152_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13065_ (.CLK(clknet_leaf_153_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13066_ (.CLK(clknet_leaf_153_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13067_ (.CLK(clknet_leaf_159_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13068_ (.CLK(clknet_leaf_157_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13069_ (.CLK(clknet_leaf_150_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13070_ (.CLK(clknet_leaf_153_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13071_ (.CLK(clknet_leaf_154_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13072_ (.CLK(clknet_leaf_154_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13073_ (.CLK(clknet_leaf_154_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13074_ (.CLK(clknet_leaf_154_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13075_ (.CLK(clknet_leaf_150_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13076_ (.CLK(clknet_leaf_149_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13077_ (.CLK(clknet_leaf_149_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13078_ (.CLK(clknet_leaf_150_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13079_ (.CLK(clknet_leaf_147_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13080_ (.CLK(clknet_leaf_146_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13081_ (.CLK(clknet_leaf_146_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13082_ (.CLK(clknet_leaf_146_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13083_ (.CLK(clknet_leaf_150_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13084_ (.CLK(clknet_leaf_150_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13085_ (.CLK(clknet_leaf_150_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13086_ (.CLK(clknet_leaf_150_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13087_ (.CLK(clknet_leaf_152_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13088_ (.CLK(clknet_leaf_151_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13089_ (.CLK(clknet_leaf_152_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13090_ (.CLK(clknet_leaf_152_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13091_ (.CLK(clknet_leaf_162_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13092_ (.CLK(clknet_leaf_163_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13093_ (.CLK(clknet_leaf_163_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13094_ (.CLK(clknet_leaf_163_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13095_ (.CLK(clknet_leaf_159_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13096_ (.CLK(clknet_leaf_159_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13097_ (.CLK(clknet_leaf_159_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13098_ (.CLK(clknet_leaf_160_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13099_ (.CLK(clknet_leaf_158_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13100_ (.CLK(clknet_leaf_160_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13101_ (.CLK(clknet_leaf_160_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13102_ (.CLK(clknet_leaf_158_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13103_ (.CLK(clknet_leaf_121_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13104_ (.CLK(clknet_leaf_121_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13105_ (.CLK(clknet_leaf_121_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13106_ (.CLK(clknet_leaf_152_clk),
    .D(net2101),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13107_ (.CLK(clknet_leaf_153_clk),
    .D(net2387),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13108_ (.CLK(clknet_leaf_153_clk),
    .D(net1914),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13109_ (.CLK(clknet_leaf_153_clk),
    .D(net2430),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13110_ (.CLK(clknet_leaf_152_clk),
    .D(net2036),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13111_ (.CLK(clknet_leaf_152_clk),
    .D(net2759),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13112_ (.CLK(clknet_leaf_153_clk),
    .D(net2397),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13113_ (.CLK(clknet_leaf_153_clk),
    .D(net1925),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13114_ (.CLK(clknet_leaf_157_clk),
    .D(net809),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13115_ (.CLK(clknet_leaf_156_clk),
    .D(net245),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13116_ (.CLK(clknet_leaf_150_clk),
    .D(net2726),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13117_ (.CLK(clknet_leaf_153_clk),
    .D(net2049),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13118_ (.CLK(clknet_leaf_154_clk),
    .D(net1789),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13119_ (.CLK(clknet_leaf_154_clk),
    .D(net1540),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13120_ (.CLK(clknet_leaf_154_clk),
    .D(net2291),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13121_ (.CLK(clknet_leaf_154_clk),
    .D(net2235),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13122_ (.CLK(clknet_leaf_151_clk),
    .D(net761),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13123_ (.CLK(clknet_leaf_149_clk),
    .D(net2308),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13124_ (.CLK(clknet_leaf_149_clk),
    .D(net1199),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13125_ (.CLK(clknet_leaf_150_clk),
    .D(net2064),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13126_ (.CLK(clknet_leaf_147_clk),
    .D(net2054),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13127_ (.CLK(clknet_leaf_146_clk),
    .D(net1941),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13128_ (.CLK(clknet_leaf_146_clk),
    .D(net1002),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13129_ (.CLK(clknet_leaf_146_clk),
    .D(net1010),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13130_ (.CLK(clknet_leaf_150_clk),
    .D(net1685),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13131_ (.CLK(clknet_leaf_150_clk),
    .D(net2108),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13132_ (.CLK(clknet_leaf_150_clk),
    .D(net1852),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13133_ (.CLK(clknet_leaf_150_clk),
    .D(net1823),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13134_ (.CLK(clknet_leaf_152_clk),
    .D(net2842),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13135_ (.CLK(clknet_leaf_151_clk),
    .D(net1038),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13136_ (.CLK(clknet_leaf_152_clk),
    .D(net1758),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13137_ (.CLK(clknet_leaf_152_clk),
    .D(net1393),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13138_ (.CLK(clknet_leaf_162_clk),
    .D(net2725),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13139_ (.CLK(clknet_leaf_162_clk),
    .D(net522),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13140_ (.CLK(clknet_leaf_162_clk),
    .D(net712),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13141_ (.CLK(clknet_leaf_162_clk),
    .D(net573),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13142_ (.CLK(clknet_leaf_164_clk),
    .D(net715),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13143_ (.CLK(clknet_leaf_160_clk),
    .D(net2059),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13144_ (.CLK(clknet_leaf_159_clk),
    .D(net1535),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13145_ (.CLK(clknet_leaf_159_clk),
    .D(net188),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13146_ (.CLK(clknet_leaf_159_clk),
    .D(net591),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13147_ (.CLK(clknet_leaf_160_clk),
    .D(net833),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13148_ (.CLK(clknet_leaf_160_clk),
    .D(net1009),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13149_ (.CLK(clknet_leaf_159_clk),
    .D(net390),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13150_ (.CLK(clknet_leaf_121_clk),
    .D(net2644),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13151_ (.CLK(clknet_leaf_121_clk),
    .D(net2475),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13152_ (.CLK(clknet_leaf_122_clk),
    .D(net767),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13153_ (.CLK(clknet_leaf_152_clk),
    .D(net1113),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13154_ (.CLK(clknet_leaf_153_clk),
    .D(net2721),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13155_ (.CLK(clknet_leaf_154_clk),
    .D(net646),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13156_ (.CLK(clknet_leaf_153_clk),
    .D(net2837),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13157_ (.CLK(clknet_leaf_152_clk),
    .D(net2103),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13158_ (.CLK(clknet_leaf_152_clk),
    .D(net2520),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13159_ (.CLK(clknet_leaf_153_clk),
    .D(net2383),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13160_ (.CLK(clknet_leaf_153_clk),
    .D(net2768),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13161_ (.CLK(clknet_leaf_160_clk),
    .D(net748),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13162_ (.CLK(clknet_leaf_157_clk),
    .D(net781),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13163_ (.CLK(clknet_leaf_150_clk),
    .D(net1310),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13164_ (.CLK(clknet_leaf_153_clk),
    .D(net1416),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13165_ (.CLK(clknet_leaf_154_clk),
    .D(net2693),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13166_ (.CLK(clknet_leaf_154_clk),
    .D(net2810),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13167_ (.CLK(clknet_leaf_154_clk),
    .D(net1568),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13168_ (.CLK(clknet_leaf_154_clk),
    .D(net2687),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13169_ (.CLK(clknet_leaf_146_clk),
    .D(net189),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13170_ (.CLK(clknet_leaf_149_clk),
    .D(net1813),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13171_ (.CLK(clknet_leaf_148_clk),
    .D(net429),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13172_ (.CLK(clknet_leaf_150_clk),
    .D(net1365),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13173_ (.CLK(clknet_leaf_147_clk),
    .D(net2516),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13174_ (.CLK(clknet_leaf_146_clk),
    .D(net1408),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13175_ (.CLK(clknet_leaf_146_clk),
    .D(net2583),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13176_ (.CLK(clknet_leaf_146_clk),
    .D(net1873),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13177_ (.CLK(clknet_leaf_150_clk),
    .D(net2570),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13178_ (.CLK(clknet_leaf_150_clk),
    .D(net1956),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13179_ (.CLK(clknet_leaf_150_clk),
    .D(net2654),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13180_ (.CLK(clknet_leaf_150_clk),
    .D(net1321),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13181_ (.CLK(clknet_leaf_151_clk),
    .D(net763),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13182_ (.CLK(clknet_leaf_151_clk),
    .D(net1881),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13183_ (.CLK(clknet_leaf_152_clk),
    .D(net2736),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13184_ (.CLK(clknet_leaf_152_clk),
    .D(net1043),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13185_ (.CLK(clknet_leaf_162_clk),
    .D(net2758),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13186_ (.CLK(clknet_leaf_162_clk),
    .D(net2454),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13187_ (.CLK(clknet_leaf_162_clk),
    .D(net2724),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13188_ (.CLK(clknet_leaf_162_clk),
    .D(net1627),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13189_ (.CLK(clknet_leaf_164_clk),
    .D(net1008),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13190_ (.CLK(clknet_leaf_161_clk),
    .D(net169),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13191_ (.CLK(clknet_leaf_160_clk),
    .D(net1771),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13192_ (.CLK(clknet_leaf_160_clk),
    .D(net2272),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13193_ (.CLK(clknet_leaf_159_clk),
    .D(net2891),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13194_ (.CLK(clknet_leaf_161_clk),
    .D(net170),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13195_ (.CLK(clknet_leaf_160_clk),
    .D(net861),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13196_ (.CLK(clknet_leaf_159_clk),
    .D(net2568),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13197_ (.CLK(clknet_leaf_121_clk),
    .D(net2376),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13198_ (.CLK(clknet_leaf_121_clk),
    .D(net1773),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13199_ (.CLK(clknet_leaf_121_clk),
    .D(net284),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13200_ (.CLK(clknet_leaf_152_clk),
    .D(net1531),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13201_ (.CLK(clknet_leaf_153_clk),
    .D(net1649),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13202_ (.CLK(clknet_leaf_153_clk),
    .D(net367),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13203_ (.CLK(clknet_leaf_153_clk),
    .D(net2024),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13204_ (.CLK(clknet_leaf_152_clk),
    .D(net2597),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13205_ (.CLK(clknet_leaf_152_clk),
    .D(net2949),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13206_ (.CLK(clknet_leaf_151_clk),
    .D(net772),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13207_ (.CLK(clknet_leaf_151_clk),
    .D(net771),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13208_ (.CLK(clknet_leaf_160_clk),
    .D(net827),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13209_ (.CLK(clknet_leaf_157_clk),
    .D(net1112),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13210_ (.CLK(clknet_leaf_150_clk),
    .D(net1848),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13211_ (.CLK(clknet_leaf_153_clk),
    .D(net1430),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13212_ (.CLK(clknet_leaf_153_clk),
    .D(net382),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13213_ (.CLK(clknet_leaf_153_clk),
    .D(net450),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13214_ (.CLK(clknet_leaf_154_clk),
    .D(net1203),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13215_ (.CLK(clknet_leaf_153_clk),
    .D(net377),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13216_ (.CLK(clknet_leaf_146_clk),
    .D(net1014),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13217_ (.CLK(clknet_leaf_148_clk),
    .D(net401),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13218_ (.CLK(clknet_leaf_148_clk),
    .D(net995),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13219_ (.CLK(clknet_leaf_150_clk),
    .D(net1274),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13220_ (.CLK(clknet_leaf_147_clk),
    .D(net1920),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13221_ (.CLK(clknet_leaf_146_clk),
    .D(net2678),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13222_ (.CLK(clknet_leaf_145_clk),
    .D(net801),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13223_ (.CLK(clknet_leaf_146_clk),
    .D(net2170),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13224_ (.CLK(clknet_leaf_150_clk),
    .D(net1035),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13225_ (.CLK(clknet_leaf_151_clk),
    .D(net758),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13226_ (.CLK(clknet_leaf_151_clk),
    .D(net755),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13227_ (.CLK(clknet_leaf_150_clk),
    .D(net1362),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13228_ (.CLK(clknet_leaf_146_clk),
    .D(net182),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13229_ (.CLK(clknet_leaf_151_clk),
    .D(net1859),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13230_ (.CLK(clknet_leaf_151_clk),
    .D(net648),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13231_ (.CLK(clknet_leaf_151_clk),
    .D(net678),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13232_ (.CLK(clknet_leaf_162_clk),
    .D(net2074),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13233_ (.CLK(clknet_leaf_162_clk),
    .D(net1237),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13234_ (.CLK(clknet_leaf_162_clk),
    .D(net1778),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13235_ (.CLK(clknet_leaf_162_clk),
    .D(net1174),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13236_ (.CLK(clknet_leaf_162_clk),
    .D(net278),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13237_ (.CLK(clknet_leaf_161_clk),
    .D(net1695),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13238_ (.CLK(clknet_leaf_160_clk),
    .D(net826),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13239_ (.CLK(clknet_leaf_160_clk),
    .D(net829),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13240_ (.CLK(clknet_leaf_160_clk),
    .D(net2928),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13241_ (.CLK(clknet_leaf_161_clk),
    .D(net2745),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13242_ (.CLK(clknet_leaf_149_clk),
    .D(net183),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13243_ (.CLK(clknet_leaf_159_clk),
    .D(net2839),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13244_ (.CLK(clknet_leaf_121_clk),
    .D(net2527),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _13245_ (.CLK(clknet_leaf_121_clk),
    .D(net1776),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _13246_ (.CLK(clknet_leaf_122_clk),
    .D(net749),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_2 _13247_ (.CLK(clknet_leaf_159_clk),
    .D(_00103_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _13248_ (.CLK(clknet_leaf_159_clk),
    .D(_00104_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13249_ (.CLK(clknet_leaf_159_clk),
    .D(_00105_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13250_ (.CLK(clknet_leaf_159_clk),
    .D(_00106_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13251_ (.CLK(clknet_leaf_159_clk),
    .D(_00107_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13252_ (.CLK(clknet_leaf_159_clk),
    .D(_00108_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13253_ (.CLK(clknet_leaf_159_clk),
    .D(_00109_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13254_ (.CLK(clknet_leaf_122_clk),
    .D(_00110_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ));
 sky130_fd_sc_hd__dfxtp_1 _13255_ (.CLK(clknet_leaf_122_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13256_ (.CLK(clknet_leaf_122_clk),
    .D(net1636),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13257_ (.CLK(clknet_leaf_122_clk),
    .D(net2325),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13258_ (.CLK(clknet_leaf_122_clk),
    .D(net1332),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13259_ (.CLK(clknet_leaf_148_clk),
    .D(_00011_),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _13260_ (.CLK(clknet_leaf_161_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13261_ (.CLK(clknet_leaf_150_clk),
    .D(net3115),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13262_ (.CLK(clknet_leaf_151_clk),
    .D(net3006),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13263_ (.CLK(clknet_leaf_151_clk),
    .D(net3044),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13264_ (.CLK(clknet_leaf_150_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13265_ (.CLK(clknet_leaf_146_clk),
    .D(net3003),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13266_ (.CLK(clknet_leaf_151_clk),
    .D(net386),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13267_ (.CLK(clknet_leaf_151_clk),
    .D(net3068),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13268_ (.CLK(clknet_leaf_161_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13269_ (.CLK(clknet_leaf_151_clk),
    .D(net3137),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13270_ (.CLK(clknet_leaf_151_clk),
    .D(net3098),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13271_ (.CLK(clknet_leaf_151_clk),
    .D(net3077),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13272_ (.CLK(clknet_leaf_161_clk),
    .D(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13273_ (.CLK(clknet_leaf_146_clk),
    .D(net3065),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13274_ (.CLK(clknet_leaf_146_clk),
    .D(net3134),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13275_ (.CLK(clknet_leaf_147_clk),
    .D(net3004),
    .Q(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13276_ (.CLK(clknet_leaf_159_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13277_ (.CLK(clknet_leaf_164_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13278_ (.CLK(clknet_leaf_158_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13279_ (.CLK(clknet_leaf_164_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13280_ (.CLK(clknet_leaf_165_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13281_ (.CLK(clknet_leaf_170_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13282_ (.CLK(clknet_leaf_170_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13283_ (.CLK(clknet_leaf_158_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13284_ (.CLK(clknet_leaf_168_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13285_ (.CLK(clknet_leaf_168_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13286_ (.CLK(clknet_leaf_168_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13287_ (.CLK(clknet_leaf_168_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13288_ (.CLK(clknet_leaf_164_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13289_ (.CLK(clknet_leaf_163_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13290_ (.CLK(clknet_leaf_164_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13291_ (.CLK(clknet_leaf_164_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13292_ (.CLK(clknet_leaf_166_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13293_ (.CLK(clknet_leaf_167_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13294_ (.CLK(clknet_leaf_167_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13295_ (.CLK(clknet_leaf_168_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13296_ (.CLK(clknet_leaf_121_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13297_ (.CLK(clknet_leaf_121_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13298_ (.CLK(clknet_leaf_121_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13299_ (.CLK(clknet_leaf_121_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13300_ (.CLK(clknet_leaf_165_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13301_ (.CLK(clknet_leaf_165_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13302_ (.CLK(clknet_leaf_165_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13303_ (.CLK(clknet_leaf_166_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13304_ (.CLK(clknet_leaf_163_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13305_ (.CLK(clknet_leaf_163_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13306_ (.CLK(clknet_leaf_163_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13307_ (.CLK(clknet_leaf_163_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13308_ (.CLK(clknet_leaf_172_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13309_ (.CLK(clknet_leaf_171_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13310_ (.CLK(clknet_leaf_171_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13311_ (.CLK(clknet_leaf_171_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13312_ (.CLK(clknet_leaf_171_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13313_ (.CLK(clknet_leaf_171_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13314_ (.CLK(clknet_leaf_170_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13315_ (.CLK(clknet_leaf_170_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13316_ (.CLK(clknet_leaf_170_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13317_ (.CLK(clknet_leaf_169_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13318_ (.CLK(clknet_leaf_170_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13319_ (.CLK(clknet_leaf_170_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13320_ (.CLK(clknet_leaf_167_clk),
    .D(net3244),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13321_ (.CLK(clknet_leaf_120_clk),
    .D(net3214),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13322_ (.CLK(clknet_leaf_167_clk),
    .D(net3306),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13323_ (.CLK(clknet_leaf_158_clk),
    .D(net651),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13324_ (.CLK(clknet_leaf_158_clk),
    .D(net119),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13325_ (.CLK(clknet_leaf_159_clk),
    .D(net343),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13326_ (.CLK(clknet_leaf_164_clk),
    .D(net935),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13327_ (.CLK(clknet_leaf_165_clk),
    .D(net1922),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13328_ (.CLK(clknet_leaf_165_clk),
    .D(net75),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13329_ (.CLK(clknet_leaf_176_clk),
    .D(net117),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13330_ (.CLK(clknet_leaf_164_clk),
    .D(net659),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13331_ (.CLK(clknet_leaf_168_clk),
    .D(net1296),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13332_ (.CLK(clknet_leaf_168_clk),
    .D(net2436),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13333_ (.CLK(clknet_leaf_169_clk),
    .D(net387),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13334_ (.CLK(clknet_leaf_169_clk),
    .D(net556),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13335_ (.CLK(clknet_leaf_163_clk),
    .D(net259),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13336_ (.CLK(clknet_leaf_163_clk),
    .D(net1403),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13337_ (.CLK(clknet_leaf_163_clk),
    .D(net261),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13338_ (.CLK(clknet_leaf_164_clk),
    .D(net1907),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13339_ (.CLK(clknet_leaf_166_clk),
    .D(net867),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13340_ (.CLK(clknet_leaf_167_clk),
    .D(net2873),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13341_ (.CLK(clknet_leaf_167_clk),
    .D(net2548),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13342_ (.CLK(clknet_leaf_167_clk),
    .D(net71),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13343_ (.CLK(clknet_leaf_121_clk),
    .D(net1650),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13344_ (.CLK(clknet_leaf_166_clk),
    .D(net845),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13345_ (.CLK(clknet_leaf_121_clk),
    .D(net2315),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13346_ (.CLK(clknet_leaf_125_clk),
    .D(net544),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13347_ (.CLK(clknet_leaf_165_clk),
    .D(net2634),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13348_ (.CLK(clknet_leaf_165_clk),
    .D(net2418),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13349_ (.CLK(clknet_leaf_165_clk),
    .D(net2498),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13350_ (.CLK(clknet_leaf_165_clk),
    .D(net223),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13351_ (.CLK(clknet_leaf_163_clk),
    .D(net1730),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13352_ (.CLK(clknet_leaf_162_clk),
    .D(net586),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13353_ (.CLK(clknet_leaf_163_clk),
    .D(net2132),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13354_ (.CLK(clknet_leaf_163_clk),
    .D(net2694),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13355_ (.CLK(clknet_leaf_171_clk),
    .D(net615),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13356_ (.CLK(clknet_leaf_171_clk),
    .D(net1349),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13357_ (.CLK(clknet_leaf_171_clk),
    .D(net2673),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13358_ (.CLK(clknet_leaf_171_clk),
    .D(net2081),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13359_ (.CLK(clknet_leaf_171_clk),
    .D(net2110),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13360_ (.CLK(clknet_leaf_171_clk),
    .D(net2509),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13361_ (.CLK(clknet_leaf_170_clk),
    .D(net2533),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13362_ (.CLK(clknet_leaf_170_clk),
    .D(net1638),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13363_ (.CLK(clknet_leaf_170_clk),
    .D(net2808),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13364_ (.CLK(clknet_leaf_169_clk),
    .D(net2761),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13365_ (.CLK(clknet_leaf_165_clk),
    .D(net69),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13366_ (.CLK(clknet_leaf_165_clk),
    .D(net81),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13367_ (.CLK(clknet_leaf_120_clk),
    .D(net528),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13368_ (.CLK(clknet_leaf_120_clk),
    .D(net2437),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13369_ (.CLK(clknet_leaf_167_clk),
    .D(net2804),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13370_ (.CLK(clknet_leaf_158_clk),
    .D(net1869),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13371_ (.CLK(clknet_leaf_164_clk),
    .D(net507),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13372_ (.CLK(clknet_leaf_159_clk),
    .D(net2347),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13373_ (.CLK(clknet_leaf_164_clk),
    .D(net2410),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13374_ (.CLK(clknet_leaf_164_clk),
    .D(net788),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13375_ (.CLK(clknet_leaf_164_clk),
    .D(net789),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13376_ (.CLK(clknet_leaf_170_clk),
    .D(net557),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13377_ (.CLK(clknet_leaf_164_clk),
    .D(net1937),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13378_ (.CLK(clknet_leaf_168_clk),
    .D(net2163),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13379_ (.CLK(clknet_leaf_168_clk),
    .D(net2316),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13380_ (.CLK(clknet_leaf_168_clk),
    .D(net612),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13381_ (.CLK(clknet_leaf_168_clk),
    .D(net595),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13382_ (.CLK(clknet_leaf_163_clk),
    .D(net1676),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13383_ (.CLK(clknet_leaf_163_clk),
    .D(net1855),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13384_ (.CLK(clknet_leaf_163_clk),
    .D(net2720),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13385_ (.CLK(clknet_leaf_164_clk),
    .D(net2819),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13386_ (.CLK(clknet_leaf_166_clk),
    .D(net1051),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13387_ (.CLK(clknet_leaf_166_clk),
    .D(net899),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13388_ (.CLK(clknet_leaf_167_clk),
    .D(net1280),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13389_ (.CLK(clknet_leaf_167_clk),
    .D(net2242),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13390_ (.CLK(clknet_leaf_122_clk),
    .D(net791),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13391_ (.CLK(clknet_leaf_121_clk),
    .D(net211),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13392_ (.CLK(clknet_leaf_166_clk),
    .D(net1219),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13393_ (.CLK(clknet_leaf_125_clk),
    .D(net2065),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13394_ (.CLK(clknet_leaf_165_clk),
    .D(net2332),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13395_ (.CLK(clknet_leaf_165_clk),
    .D(net1355),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13396_ (.CLK(clknet_leaf_165_clk),
    .D(net1441),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13397_ (.CLK(clknet_leaf_165_clk),
    .D(net1870),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13398_ (.CLK(clknet_leaf_163_clk),
    .D(net2346),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13399_ (.CLK(clknet_leaf_162_clk),
    .D(net2777),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13400_ (.CLK(clknet_leaf_162_clk),
    .D(net754),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13401_ (.CLK(clknet_leaf_163_clk),
    .D(net2190),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13402_ (.CLK(clknet_leaf_171_clk),
    .D(net1623),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13403_ (.CLK(clknet_leaf_171_clk),
    .D(net2137),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13404_ (.CLK(clknet_leaf_171_clk),
    .D(net2086),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13405_ (.CLK(clknet_leaf_171_clk),
    .D(net1987),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13406_ (.CLK(clknet_leaf_171_clk),
    .D(net2419),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13407_ (.CLK(clknet_leaf_171_clk),
    .D(net1542),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13408_ (.CLK(clknet_leaf_170_clk),
    .D(net1847),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13409_ (.CLK(clknet_leaf_170_clk),
    .D(net1170),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13410_ (.CLK(clknet_leaf_170_clk),
    .D(net1528),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13411_ (.CLK(clknet_leaf_169_clk),
    .D(net1679),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13412_ (.CLK(clknet_leaf_165_clk),
    .D(net1368),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13413_ (.CLK(clknet_leaf_170_clk),
    .D(net122),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13414_ (.CLK(clknet_leaf_167_clk),
    .D(net516),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13415_ (.CLK(clknet_leaf_120_clk),
    .D(net2015),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13416_ (.CLK(clknet_leaf_167_clk),
    .D(net1846),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13417_ (.CLK(clknet_leaf_159_clk),
    .D(net453),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13418_ (.CLK(clknet_leaf_164_clk),
    .D(net1375),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13419_ (.CLK(clknet_leaf_159_clk),
    .D(net2609),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13420_ (.CLK(clknet_leaf_164_clk),
    .D(net1005),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13421_ (.CLK(clknet_leaf_164_clk),
    .D(net1157),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13422_ (.CLK(clknet_leaf_164_clk),
    .D(net2298),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13423_ (.CLK(clknet_leaf_164_clk),
    .D(net79),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13424_ (.CLK(clknet_leaf_158_clk),
    .D(net116),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13425_ (.CLK(clknet_leaf_168_clk),
    .D(net1916),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13426_ (.CLK(clknet_leaf_168_clk),
    .D(net2541),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13427_ (.CLK(clknet_leaf_168_clk),
    .D(net1411),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13428_ (.CLK(clknet_leaf_168_clk),
    .D(net2464),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13429_ (.CLK(clknet_leaf_163_clk),
    .D(net2511),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13430_ (.CLK(clknet_leaf_162_clk),
    .D(net711),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13431_ (.CLK(clknet_leaf_163_clk),
    .D(net2543),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13432_ (.CLK(clknet_leaf_164_clk),
    .D(net1824),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13433_ (.CLK(clknet_leaf_166_clk),
    .D(net900),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13434_ (.CLK(clknet_leaf_166_clk),
    .D(net868),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13435_ (.CLK(clknet_leaf_167_clk),
    .D(net2020),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13436_ (.CLK(clknet_leaf_167_clk),
    .D(net2824),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13437_ (.CLK(clknet_leaf_125_clk),
    .D(net289),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13438_ (.CLK(clknet_leaf_121_clk),
    .D(net2032),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13439_ (.CLK(clknet_leaf_121_clk),
    .D(net226),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13440_ (.CLK(clknet_leaf_125_clk),
    .D(net2750),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13441_ (.CLK(clknet_leaf_165_clk),
    .D(net1109),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13442_ (.CLK(clknet_leaf_165_clk),
    .D(net1729),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13443_ (.CLK(clknet_leaf_165_clk),
    .D(net2786),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13444_ (.CLK(clknet_leaf_165_clk),
    .D(net1641),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13445_ (.CLK(clknet_leaf_125_clk),
    .D(net653),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13446_ (.CLK(clknet_leaf_162_clk),
    .D(net2403),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13447_ (.CLK(clknet_leaf_162_clk),
    .D(net2539),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13448_ (.CLK(clknet_leaf_162_clk),
    .D(net743),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13449_ (.CLK(clknet_leaf_171_clk),
    .D(net2002),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13450_ (.CLK(clknet_leaf_170_clk),
    .D(net597),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13451_ (.CLK(clknet_leaf_170_clk),
    .D(net690),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13452_ (.CLK(clknet_leaf_171_clk),
    .D(net1894),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13453_ (.CLK(clknet_leaf_171_clk),
    .D(net1253),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13454_ (.CLK(clknet_leaf_171_clk),
    .D(net1347),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13455_ (.CLK(clknet_leaf_170_clk),
    .D(net2297),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13456_ (.CLK(clknet_leaf_170_clk),
    .D(net2145),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13457_ (.CLK(clknet_leaf_170_clk),
    .D(net2127),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13458_ (.CLK(clknet_leaf_170_clk),
    .D(net704),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13459_ (.CLK(clknet_leaf_165_clk),
    .D(net2544),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13460_ (.CLK(clknet_leaf_165_clk),
    .D(net70),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13461_ (.CLK(clknet_leaf_120_clk),
    .D(net527),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _13462_ (.CLK(clknet_leaf_120_clk),
    .D(net2394),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _13463_ (.CLK(clknet_leaf_167_clk),
    .D(net1985),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _13464_ (.CLK(clknet_leaf_169_clk),
    .D(_00111_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _13465_ (.CLK(clknet_leaf_169_clk),
    .D(_00112_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13466_ (.CLK(clknet_leaf_169_clk),
    .D(_00113_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13467_ (.CLK(clknet_leaf_169_clk),
    .D(_00114_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13468_ (.CLK(clknet_leaf_169_clk),
    .D(_00115_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13469_ (.CLK(clknet_leaf_169_clk),
    .D(_00116_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13470_ (.CLK(clknet_leaf_169_clk),
    .D(_00117_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13471_ (.CLK(clknet_leaf_24_clk),
    .D(_00118_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ));
 sky130_fd_sc_hd__dfxtp_1 _13472_ (.CLK(clknet_leaf_168_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13473_ (.CLK(clknet_leaf_168_clk),
    .D(net2620),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13474_ (.CLK(clknet_leaf_167_clk),
    .D(net78),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13475_ (.CLK(clknet_leaf_167_clk),
    .D(net1882),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13476_ (.CLK(clknet_leaf_158_clk),
    .D(_00004_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _13477_ (.CLK(clknet_leaf_163_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13478_ (.CLK(clknet_leaf_163_clk),
    .D(net3062),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13479_ (.CLK(clknet_leaf_166_clk),
    .D(net3021),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13480_ (.CLK(clknet_leaf_166_clk),
    .D(net3051),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13481_ (.CLK(clknet_leaf_163_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13482_ (.CLK(clknet_leaf_166_clk),
    .D(net3038),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13483_ (.CLK(clknet_leaf_166_clk),
    .D(net3022),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13484_ (.CLK(clknet_leaf_163_clk),
    .D(net2956),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13485_ (.CLK(clknet_leaf_170_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13486_ (.CLK(clknet_leaf_166_clk),
    .D(net270),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13487_ (.CLK(clknet_leaf_165_clk),
    .D(net2951),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13488_ (.CLK(clknet_leaf_165_clk),
    .D(net3040),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13489_ (.CLK(clknet_leaf_170_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13490_ (.CLK(clknet_leaf_166_clk),
    .D(net750),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13491_ (.CLK(clknet_leaf_166_clk),
    .D(net3130),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13492_ (.CLK(clknet_leaf_166_clk),
    .D(net3104),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13493_ (.CLK(clknet_leaf_155_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13494_ (.CLK(clknet_leaf_155_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13495_ (.CLK(clknet_leaf_155_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13496_ (.CLK(clknet_leaf_155_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13497_ (.CLK(clknet_leaf_155_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13498_ (.CLK(clknet_leaf_179_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13499_ (.CLK(clknet_leaf_156_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13500_ (.CLK(clknet_leaf_155_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13501_ (.CLK(clknet_leaf_157_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13502_ (.CLK(clknet_leaf_157_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13503_ (.CLK(clknet_leaf_157_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13504_ (.CLK(clknet_leaf_157_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13505_ (.CLK(clknet_leaf_156_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13506_ (.CLK(clknet_leaf_156_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13507_ (.CLK(clknet_leaf_156_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13508_ (.CLK(clknet_leaf_156_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13509_ (.CLK(clknet_leaf_179_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13510_ (.CLK(clknet_leaf_179_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13511_ (.CLK(clknet_leaf_177_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13512_ (.CLK(clknet_leaf_178_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13513_ (.CLK(clknet_leaf_181_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13514_ (.CLK(clknet_leaf_180_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13515_ (.CLK(clknet_leaf_180_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13516_ (.CLK(clknet_leaf_180_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13517_ (.CLK(clknet_leaf_178_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13518_ (.CLK(clknet_leaf_178_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13519_ (.CLK(clknet_leaf_178_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13520_ (.CLK(clknet_leaf_178_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13521_ (.CLK(clknet_leaf_181_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13522_ (.CLK(clknet_leaf_180_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13523_ (.CLK(clknet_leaf_180_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13524_ (.CLK(clknet_leaf_180_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13525_ (.CLK(clknet_leaf_176_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13526_ (.CLK(clknet_leaf_175_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13527_ (.CLK(clknet_leaf_176_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13528_ (.CLK(clknet_leaf_176_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13529_ (.CLK(clknet_leaf_158_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13530_ (.CLK(clknet_leaf_158_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13531_ (.CLK(clknet_leaf_176_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13532_ (.CLK(clknet_leaf_158_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13533_ (.CLK(clknet_leaf_177_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13534_ (.CLK(clknet_leaf_175_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13535_ (.CLK(clknet_leaf_177_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13536_ (.CLK(clknet_leaf_177_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13537_ (.CLK(clknet_leaf_120_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13538_ (.CLK(clknet_leaf_120_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13539_ (.CLK(clknet_leaf_120_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13540_ (.CLK(clknet_leaf_155_clk),
    .D(net2318),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13541_ (.CLK(clknet_leaf_155_clk),
    .D(net1272),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13542_ (.CLK(clknet_leaf_155_clk),
    .D(net1794),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13543_ (.CLK(clknet_leaf_154_clk),
    .D(net488),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13544_ (.CLK(clknet_leaf_155_clk),
    .D(net1958),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13545_ (.CLK(clknet_leaf_155_clk),
    .D(net65),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13546_ (.CLK(clknet_leaf_154_clk),
    .D(net551),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13547_ (.CLK(clknet_leaf_155_clk),
    .D(net1184),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13548_ (.CLK(clknet_leaf_157_clk),
    .D(net894),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13549_ (.CLK(clknet_leaf_157_clk),
    .D(net1121),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13550_ (.CLK(clknet_leaf_157_clk),
    .D(net949),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13551_ (.CLK(clknet_leaf_157_clk),
    .D(net1122),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13552_ (.CLK(clknet_leaf_156_clk),
    .D(net2739),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13553_ (.CLK(clknet_leaf_156_clk),
    .D(net2594),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13554_ (.CLK(clknet_leaf_156_clk),
    .D(net2051),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13555_ (.CLK(clknet_leaf_156_clk),
    .D(net2888),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13556_ (.CLK(clknet_leaf_179_clk),
    .D(net828),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13557_ (.CLK(clknet_leaf_156_clk),
    .D(net62),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13558_ (.CLK(clknet_leaf_177_clk),
    .D(net1893),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13559_ (.CLK(clknet_leaf_177_clk),
    .D(net619),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13560_ (.CLK(clknet_leaf_181_clk),
    .D(net2427),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13561_ (.CLK(clknet_leaf_180_clk),
    .D(net1827),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13562_ (.CLK(clknet_leaf_180_clk),
    .D(net2129),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13563_ (.CLK(clknet_leaf_180_clk),
    .D(net2535),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13564_ (.CLK(clknet_leaf_178_clk),
    .D(net1890),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13565_ (.CLK(clknet_leaf_178_clk),
    .D(net2651),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13566_ (.CLK(clknet_leaf_177_clk),
    .D(net571),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13567_ (.CLK(clknet_leaf_178_clk),
    .D(net1305),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13568_ (.CLK(clknet_leaf_181_clk),
    .D(net2886),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13569_ (.CLK(clknet_leaf_180_clk),
    .D(net2795),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13570_ (.CLK(clknet_leaf_180_clk),
    .D(net2481),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13571_ (.CLK(clknet_leaf_180_clk),
    .D(net2580),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13572_ (.CLK(clknet_leaf_175_clk),
    .D(net304),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13573_ (.CLK(clknet_leaf_175_clk),
    .D(net2273),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13574_ (.CLK(clknet_leaf_176_clk),
    .D(net1050),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13575_ (.CLK(clknet_leaf_176_clk),
    .D(net2662),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13576_ (.CLK(clknet_leaf_158_clk),
    .D(net1213),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13577_ (.CLK(clknet_leaf_158_clk),
    .D(net2933),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13578_ (.CLK(clknet_leaf_176_clk),
    .D(net1779),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13579_ (.CLK(clknet_leaf_177_clk),
    .D(net95),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13580_ (.CLK(clknet_leaf_177_clk),
    .D(net1397),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13581_ (.CLK(clknet_leaf_175_clk),
    .D(net2351),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13582_ (.CLK(clknet_leaf_177_clk),
    .D(net1537),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13583_ (.CLK(clknet_leaf_175_clk),
    .D(net412),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13584_ (.CLK(clknet_leaf_119_clk),
    .D(net111),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13585_ (.CLK(clknet_leaf_120_clk),
    .D(net2039),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13586_ (.CLK(clknet_leaf_120_clk),
    .D(net2715),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13587_ (.CLK(clknet_leaf_155_clk),
    .D(net2378),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13588_ (.CLK(clknet_leaf_155_clk),
    .D(net2261),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13589_ (.CLK(clknet_leaf_154_clk),
    .D(net459),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13590_ (.CLK(clknet_leaf_155_clk),
    .D(net449),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13591_ (.CLK(clknet_leaf_155_clk),
    .D(net2598),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13592_ (.CLK(clknet_leaf_155_clk),
    .D(net2204),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13593_ (.CLK(clknet_leaf_154_clk),
    .D(net2661),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13594_ (.CLK(clknet_leaf_155_clk),
    .D(net2171),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13595_ (.CLK(clknet_leaf_157_clk),
    .D(net1495),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13596_ (.CLK(clknet_leaf_156_clk),
    .D(net241),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13597_ (.CLK(clknet_leaf_156_clk),
    .D(net251),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13598_ (.CLK(clknet_leaf_157_clk),
    .D(net1673),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13599_ (.CLK(clknet_leaf_156_clk),
    .D(net2627),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13600_ (.CLK(clknet_leaf_156_clk),
    .D(net1763),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13601_ (.CLK(clknet_leaf_154_clk),
    .D(net513),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13602_ (.CLK(clknet_leaf_156_clk),
    .D(net2299),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13603_ (.CLK(clknet_leaf_156_clk),
    .D(net60),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13604_ (.CLK(clknet_leaf_156_clk),
    .D(net2529),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13605_ (.CLK(clknet_leaf_177_clk),
    .D(net1967),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13606_ (.CLK(clknet_leaf_177_clk),
    .D(net1549),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13607_ (.CLK(clknet_leaf_181_clk),
    .D(net2717),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13608_ (.CLK(clknet_leaf_179_clk),
    .D(net2889),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13609_ (.CLK(clknet_leaf_179_clk),
    .D(net2915),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13610_ (.CLK(clknet_leaf_180_clk),
    .D(net2323),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13611_ (.CLK(clknet_leaf_178_clk),
    .D(net2755),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13612_ (.CLK(clknet_leaf_178_clk),
    .D(net1312),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13613_ (.CLK(clknet_leaf_177_clk),
    .D(net2189),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13614_ (.CLK(clknet_leaf_178_clk),
    .D(net1795),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13615_ (.CLK(clknet_leaf_181_clk),
    .D(net2895),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13616_ (.CLK(clknet_leaf_180_clk),
    .D(net2120),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13617_ (.CLK(clknet_leaf_180_clk),
    .D(net1422),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13618_ (.CLK(clknet_leaf_180_clk),
    .D(net2262),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13619_ (.CLK(clknet_leaf_176_clk),
    .D(net737),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13620_ (.CLK(clknet_leaf_175_clk),
    .D(net1571),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13621_ (.CLK(clknet_leaf_176_clk),
    .D(net1439),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13622_ (.CLK(clknet_leaf_176_clk),
    .D(net1095),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13623_ (.CLK(clknet_leaf_158_clk),
    .D(net2201),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13624_ (.CLK(clknet_leaf_158_clk),
    .D(net2307),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13625_ (.CLK(clknet_leaf_176_clk),
    .D(net1153),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13626_ (.CLK(clknet_leaf_158_clk),
    .D(net85),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13627_ (.CLK(clknet_leaf_177_clk),
    .D(net2083),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13628_ (.CLK(clknet_leaf_176_clk),
    .D(net752),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13629_ (.CLK(clknet_leaf_177_clk),
    .D(net2350),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13630_ (.CLK(clknet_leaf_177_clk),
    .D(net680),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13631_ (.CLK(clknet_leaf_119_clk),
    .D(net2615),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13632_ (.CLK(clknet_leaf_119_clk),
    .D(net104),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13633_ (.CLK(clknet_leaf_120_clk),
    .D(net2885),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13634_ (.CLK(clknet_leaf_155_clk),
    .D(net2487),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13635_ (.CLK(clknet_leaf_155_clk),
    .D(net2870),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13636_ (.CLK(clknet_leaf_154_clk),
    .D(net1697),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13637_ (.CLK(clknet_leaf_154_clk),
    .D(net534),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13638_ (.CLK(clknet_leaf_155_clk),
    .D(net2645),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13639_ (.CLK(clknet_leaf_155_clk),
    .D(net1919),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13640_ (.CLK(clknet_leaf_154_clk),
    .D(net1980),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13641_ (.CLK(clknet_leaf_154_clk),
    .D(net582),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13642_ (.CLK(clknet_leaf_159_clk),
    .D(net234),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13643_ (.CLK(clknet_leaf_156_clk),
    .D(net2545),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13644_ (.CLK(clknet_leaf_157_clk),
    .D(net844),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13645_ (.CLK(clknet_leaf_157_clk),
    .D(net2499),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13646_ (.CLK(clknet_leaf_153_clk),
    .D(net554),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13647_ (.CLK(clknet_leaf_156_clk),
    .D(net1402),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13648_ (.CLK(clknet_leaf_154_clk),
    .D(net2334),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13649_ (.CLK(clknet_leaf_156_clk),
    .D(net2070),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13650_ (.CLK(clknet_leaf_156_clk),
    .D(net1462),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13651_ (.CLK(clknet_leaf_156_clk),
    .D(net1787),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13652_ (.CLK(clknet_leaf_157_clk),
    .D(net99),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13653_ (.CLK(clknet_leaf_177_clk),
    .D(net1478),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13654_ (.CLK(clknet_leaf_181_clk),
    .D(net1134),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13655_ (.CLK(clknet_leaf_179_clk),
    .D(net822),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13656_ (.CLK(clknet_leaf_179_clk),
    .D(net830),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13657_ (.CLK(clknet_leaf_155_clk),
    .D(net87),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13658_ (.CLK(clknet_leaf_178_clk),
    .D(net1098),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13659_ (.CLK(clknet_leaf_178_clk),
    .D(net2181),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13660_ (.CLK(clknet_leaf_177_clk),
    .D(net1198),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13661_ (.CLK(clknet_leaf_177_clk),
    .D(net485),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13662_ (.CLK(clknet_leaf_181_clk),
    .D(net973),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13663_ (.CLK(clknet_leaf_180_clk),
    .D(net2774),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13664_ (.CLK(clknet_leaf_180_clk),
    .D(net1617),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13665_ (.CLK(clknet_leaf_180_clk),
    .D(net2478),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13666_ (.CLK(clknet_leaf_176_clk),
    .D(net1560),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13667_ (.CLK(clknet_leaf_176_clk),
    .D(net768),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13668_ (.CLK(clknet_leaf_176_clk),
    .D(net1955),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13669_ (.CLK(clknet_leaf_176_clk),
    .D(net1181),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13670_ (.CLK(clknet_leaf_158_clk),
    .D(net2683),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13671_ (.CLK(clknet_leaf_158_clk),
    .D(net2305),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13672_ (.CLK(clknet_leaf_158_clk),
    .D(net80),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13673_ (.CLK(clknet_leaf_158_clk),
    .D(net1703),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13674_ (.CLK(clknet_leaf_177_clk),
    .D(net1507),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13675_ (.CLK(clknet_leaf_176_clk),
    .D(net941),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13676_ (.CLK(clknet_leaf_177_clk),
    .D(net1320),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13677_ (.CLK(clknet_leaf_177_clk),
    .D(net2048),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13678_ (.CLK(clknet_leaf_119_clk),
    .D(net2836),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _13679_ (.CLK(clknet_leaf_119_clk),
    .D(net2380),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _13680_ (.CLK(clknet_leaf_120_clk),
    .D(net2924),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _13681_ (.CLK(clknet_leaf_158_clk),
    .D(_00119_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _13682_ (.CLK(clknet_leaf_159_clk),
    .D(_00120_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13683_ (.CLK(clknet_leaf_157_clk),
    .D(_00121_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13684_ (.CLK(clknet_leaf_157_clk),
    .D(_00122_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13685_ (.CLK(clknet_leaf_158_clk),
    .D(_00123_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13686_ (.CLK(clknet_leaf_158_clk),
    .D(_00124_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13687_ (.CLK(clknet_leaf_158_clk),
    .D(_00125_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13688_ (.CLK(clknet_leaf_68_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13689_ (.CLK(clknet_leaf_68_clk),
    .D(net1180),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13690_ (.CLK(clknet_leaf_69_clk),
    .D(net57),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13691_ (.CLK(clknet_leaf_69_clk),
    .D(net2078),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13692_ (.CLK(clknet_leaf_157_clk),
    .D(_00005_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _13693_ (.CLK(clknet_leaf_176_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13694_ (.CLK(clknet_leaf_178_clk),
    .D(net3000),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13695_ (.CLK(clknet_leaf_178_clk),
    .D(net3064),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13696_ (.CLK(clknet_leaf_178_clk),
    .D(net3061),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13697_ (.CLK(clknet_leaf_178_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13698_ (.CLK(clknet_leaf_178_clk),
    .D(net3093),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13699_ (.CLK(clknet_leaf_178_clk),
    .D(net3071),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13700_ (.CLK(clknet_leaf_178_clk),
    .D(net3092),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13701_ (.CLK(clknet_leaf_177_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13702_ (.CLK(clknet_leaf_179_clk),
    .D(net3128),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13703_ (.CLK(clknet_leaf_179_clk),
    .D(net3013),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13704_ (.CLK(clknet_leaf_179_clk),
    .D(net3039),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13705_ (.CLK(clknet_leaf_177_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13706_ (.CLK(clknet_leaf_179_clk),
    .D(net3139),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13707_ (.CLK(clknet_leaf_156_clk),
    .D(net157),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13708_ (.CLK(clknet_leaf_156_clk),
    .D(net3111),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13709_ (.CLK(clknet_leaf_182_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13710_ (.CLK(clknet_leaf_181_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13711_ (.CLK(clknet_leaf_182_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13712_ (.CLK(clknet_leaf_181_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13713_ (.CLK(clknet_leaf_183_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13714_ (.CLK(clknet_leaf_183_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13715_ (.CLK(clknet_leaf_183_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13716_ (.CLK(clknet_leaf_183_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13717_ (.CLK(clknet_leaf_175_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13718_ (.CLK(clknet_leaf_181_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13719_ (.CLK(clknet_leaf_178_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13720_ (.CLK(clknet_leaf_185_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13721_ (.CLK(clknet_leaf_182_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13722_ (.CLK(clknet_leaf_182_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13723_ (.CLK(clknet_leaf_182_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13724_ (.CLK(clknet_leaf_183_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13725_ (.CLK(clknet_leaf_185_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13726_ (.CLK(clknet_leaf_185_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13727_ (.CLK(clknet_leaf_184_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13728_ (.CLK(clknet_leaf_185_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13729_ (.CLK(clknet_leaf_188_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13730_ (.CLK(clknet_leaf_189_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13731_ (.CLK(clknet_leaf_184_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13732_ (.CLK(clknet_leaf_189_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13733_ (.CLK(clknet_leaf_188_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13734_ (.CLK(clknet_leaf_185_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13735_ (.CLK(clknet_leaf_184_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13736_ (.CLK(clknet_leaf_185_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13737_ (.CLK(clknet_leaf_189_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13738_ (.CLK(clknet_leaf_188_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13739_ (.CLK(clknet_leaf_188_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13740_ (.CLK(clknet_leaf_190_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13741_ (.CLK(clknet_leaf_173_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13742_ (.CLK(clknet_leaf_174_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13743_ (.CLK(clknet_leaf_174_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13744_ (.CLK(clknet_leaf_174_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13745_ (.CLK(clknet_leaf_173_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13746_ (.CLK(clknet_leaf_175_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13747_ (.CLK(clknet_leaf_174_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13748_ (.CLK(clknet_leaf_174_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13749_ (.CLK(clknet_leaf_185_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13750_ (.CLK(clknet_leaf_185_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13751_ (.CLK(clknet_leaf_185_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13752_ (.CLK(clknet_leaf_185_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13753_ (.CLK(clknet_leaf_69_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13754_ (.CLK(clknet_leaf_69_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13755_ (.CLK(clknet_leaf_69_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13756_ (.CLK(clknet_leaf_181_clk),
    .D(net434),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13757_ (.CLK(clknet_leaf_181_clk),
    .D(net1533),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13758_ (.CLK(clknet_leaf_182_clk),
    .D(net2572),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13759_ (.CLK(clknet_leaf_181_clk),
    .D(net2448),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13760_ (.CLK(clknet_leaf_183_clk),
    .D(net1493),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13761_ (.CLK(clknet_leaf_182_clk),
    .D(net661),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13762_ (.CLK(clknet_leaf_183_clk),
    .D(net2611),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13763_ (.CLK(clknet_leaf_183_clk),
    .D(net2681),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13764_ (.CLK(clknet_leaf_175_clk),
    .D(net2621),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13765_ (.CLK(clknet_leaf_181_clk),
    .D(net2013),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13766_ (.CLK(clknet_leaf_178_clk),
    .D(net1810),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13767_ (.CLK(clknet_leaf_185_clk),
    .D(net1352),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13768_ (.CLK(clknet_leaf_182_clk),
    .D(net2599),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13769_ (.CLK(clknet_leaf_181_clk),
    .D(net504),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13770_ (.CLK(clknet_leaf_183_clk),
    .D(net394),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13771_ (.CLK(clknet_leaf_183_clk),
    .D(net2156),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13772_ (.CLK(clknet_leaf_182_clk),
    .D(net677),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13773_ (.CLK(clknet_leaf_182_clk),
    .D(net742),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13774_ (.CLK(clknet_leaf_186_clk),
    .D(net190),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13775_ (.CLK(clknet_leaf_185_clk),
    .D(net2404),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13776_ (.CLK(clknet_leaf_189_clk),
    .D(net82),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13777_ (.CLK(clknet_leaf_189_clk),
    .D(net1548),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13778_ (.CLK(clknet_leaf_183_clk),
    .D(net198),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13779_ (.CLK(clknet_leaf_183_clk),
    .D(net760),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13780_ (.CLK(clknet_leaf_188_clk),
    .D(net2080),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13781_ (.CLK(clknet_leaf_182_clk),
    .D(net594),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13782_ (.CLK(clknet_leaf_184_clk),
    .D(net1242),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13783_ (.CLK(clknet_leaf_185_clk),
    .D(net2796),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13784_ (.CLK(clknet_leaf_189_clk),
    .D(net1726),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13785_ (.CLK(clknet_leaf_189_clk),
    .D(net73),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13786_ (.CLK(clknet_leaf_188_clk),
    .D(net2872),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13787_ (.CLK(clknet_leaf_190_clk),
    .D(net1498),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13788_ (.CLK(clknet_leaf_173_clk),
    .D(net2133),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13789_ (.CLK(clknet_leaf_174_clk),
    .D(net2445),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13790_ (.CLK(clknet_leaf_174_clk),
    .D(net987),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13791_ (.CLK(clknet_leaf_173_clk),
    .D(net345),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13792_ (.CLK(clknet_leaf_174_clk),
    .D(net150),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13793_ (.CLK(clknet_leaf_174_clk),
    .D(net779),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13794_ (.CLK(clknet_leaf_173_clk),
    .D(net457),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13795_ (.CLK(clknet_leaf_174_clk),
    .D(net1651),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13796_ (.CLK(clknet_leaf_186_clk),
    .D(net671),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13797_ (.CLK(clknet_leaf_175_clk),
    .D(net424),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13798_ (.CLK(clknet_leaf_185_clk),
    .D(net2659),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13799_ (.CLK(clknet_leaf_174_clk),
    .D(net799),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13800_ (.CLK(clknet_leaf_69_clk),
    .D(net2875),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13801_ (.CLK(clknet_leaf_69_clk),
    .D(net1668),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13802_ (.CLK(clknet_leaf_69_clk),
    .D(net1405),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13803_ (.CLK(clknet_leaf_181_clk),
    .D(net1690),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13804_ (.CLK(clknet_leaf_180_clk),
    .D(net348),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13805_ (.CLK(clknet_leaf_182_clk),
    .D(net2794),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13806_ (.CLK(clknet_leaf_181_clk),
    .D(net2803),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13807_ (.CLK(clknet_leaf_183_clk),
    .D(net2218),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13808_ (.CLK(clknet_leaf_183_clk),
    .D(net514),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13809_ (.CLK(clknet_leaf_183_clk),
    .D(net2016),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13810_ (.CLK(clknet_leaf_183_clk),
    .D(net1414),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13811_ (.CLK(clknet_leaf_175_clk),
    .D(net1489),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13812_ (.CLK(clknet_leaf_181_clk),
    .D(net2883),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13813_ (.CLK(clknet_leaf_181_clk),
    .D(net722),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13814_ (.CLK(clknet_leaf_185_clk),
    .D(net2354),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13815_ (.CLK(clknet_leaf_182_clk),
    .D(net2444),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13816_ (.CLK(clknet_leaf_181_clk),
    .D(net2595),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13817_ (.CLK(clknet_leaf_182_clk),
    .D(net451),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13818_ (.CLK(clknet_leaf_182_clk),
    .D(net536),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13819_ (.CLK(clknet_leaf_181_clk),
    .D(net564),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13820_ (.CLK(clknet_leaf_182_clk),
    .D(net2618),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13821_ (.CLK(clknet_leaf_186_clk),
    .D(net1148),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13822_ (.CLK(clknet_leaf_185_clk),
    .D(net1499),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13823_ (.CLK(clknet_leaf_189_clk),
    .D(net1000),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13824_ (.CLK(clknet_leaf_189_clk),
    .D(net837),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13825_ (.CLK(clknet_leaf_184_clk),
    .D(net2413),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13826_ (.CLK(clknet_leaf_189_clk),
    .D(net74),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13827_ (.CLK(clknet_leaf_188_clk),
    .D(net1400),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13828_ (.CLK(clknet_leaf_182_clk),
    .D(net1621),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13829_ (.CLK(clknet_leaf_184_clk),
    .D(net858),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13830_ (.CLK(clknet_leaf_185_clk),
    .D(net2729),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13831_ (.CLK(clknet_leaf_189_clk),
    .D(net895),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13832_ (.CLK(clknet_leaf_188_clk),
    .D(net3100),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13833_ (.CLK(clknet_leaf_188_clk),
    .D(net2680),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13834_ (.CLK(clknet_leaf_187_clk),
    .D(net478),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13835_ (.CLK(clknet_leaf_173_clk),
    .D(net1952),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13836_ (.CLK(clknet_leaf_175_clk),
    .D(net244),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13837_ (.CLK(clknet_leaf_176_clk),
    .D(net325),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13838_ (.CLK(clknet_leaf_173_clk),
    .D(net1947),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13839_ (.CLK(clknet_leaf_173_clk),
    .D(net301),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13840_ (.CLK(clknet_leaf_175_clk),
    .D(net246),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13841_ (.CLK(clknet_leaf_173_clk),
    .D(net2695),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13842_ (.CLK(clknet_leaf_174_clk),
    .D(net1100),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13843_ (.CLK(clknet_leaf_185_clk),
    .D(net430),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13844_ (.CLK(clknet_leaf_175_clk),
    .D(net2282),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13845_ (.CLK(clknet_leaf_185_clk),
    .D(net2317),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13846_ (.CLK(clknet_leaf_174_clk),
    .D(net2012),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13847_ (.CLK(clknet_leaf_69_clk),
    .D(net2641),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13848_ (.CLK(clknet_leaf_69_clk),
    .D(net1333),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13849_ (.CLK(clknet_leaf_120_clk),
    .D(net155),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13850_ (.CLK(clknet_leaf_180_clk),
    .D(net362),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13851_ (.CLK(clknet_leaf_180_clk),
    .D(net2462),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13852_ (.CLK(clknet_leaf_181_clk),
    .D(net685),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13853_ (.CLK(clknet_leaf_181_clk),
    .D(net1736),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13854_ (.CLK(clknet_leaf_183_clk),
    .D(net1466),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13855_ (.CLK(clknet_leaf_182_clk),
    .D(net660),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13856_ (.CLK(clknet_leaf_183_clk),
    .D(net2806),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13857_ (.CLK(clknet_leaf_183_clk),
    .D(net2571),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13858_ (.CLK(clknet_leaf_178_clk),
    .D(net469),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13859_ (.CLK(clknet_leaf_178_clk),
    .D(net460),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13860_ (.CLK(clknet_leaf_178_clk),
    .D(net369),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13861_ (.CLK(clknet_leaf_185_clk),
    .D(net1377),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13862_ (.CLK(clknet_leaf_182_clk),
    .D(net1817),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13863_ (.CLK(clknet_leaf_180_clk),
    .D(net524),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13864_ (.CLK(clknet_leaf_182_clk),
    .D(net2322),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13865_ (.CLK(clknet_leaf_182_clk),
    .D(net2312),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13866_ (.CLK(clknet_leaf_182_clk),
    .D(net610),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13867_ (.CLK(clknet_leaf_182_clk),
    .D(net2760),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13868_ (.CLK(clknet_leaf_184_clk),
    .D(net1428),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13869_ (.CLK(clknet_leaf_185_clk),
    .D(net2042),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13870_ (.CLK(clknet_leaf_189_clk),
    .D(net831),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13871_ (.CLK(clknet_leaf_189_clk),
    .D(net989),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13872_ (.CLK(clknet_leaf_184_clk),
    .D(net903),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13873_ (.CLK(clknet_leaf_183_clk),
    .D(net617),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13874_ (.CLK(clknet_leaf_188_clk),
    .D(net1090),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13875_ (.CLK(clknet_leaf_181_clk),
    .D(net468),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13876_ (.CLK(clknet_leaf_184_clk),
    .D(net918),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13877_ (.CLK(clknet_leaf_185_clk),
    .D(net2213),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13878_ (.CLK(clknet_leaf_188_clk),
    .D(net3091),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13879_ (.CLK(clknet_leaf_188_clk),
    .D(net1839),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13880_ (.CLK(clknet_leaf_188_clk),
    .D(net2017),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13881_ (.CLK(clknet_leaf_187_clk),
    .D(net1360),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13882_ (.CLK(clknet_leaf_171_clk),
    .D(net652),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13883_ (.CLK(clknet_leaf_175_clk),
    .D(net1866),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13884_ (.CLK(clknet_leaf_176_clk),
    .D(net1381),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13885_ (.CLK(clknet_leaf_174_clk),
    .D(net138),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13886_ (.CLK(clknet_leaf_173_clk),
    .D(net2224),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13887_ (.CLK(clknet_leaf_174_clk),
    .D(net790),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13888_ (.CLK(clknet_leaf_174_clk),
    .D(net132),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13889_ (.CLK(clknet_leaf_174_clk),
    .D(net1056),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13890_ (.CLK(clknet_leaf_185_clk),
    .D(net2447),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13891_ (.CLK(clknet_leaf_175_clk),
    .D(net1951),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13892_ (.CLK(clknet_leaf_185_clk),
    .D(net2619),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13893_ (.CLK(clknet_leaf_174_clk),
    .D(net905),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13894_ (.CLK(clknet_leaf_69_clk),
    .D(net1814),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _13895_ (.CLK(clknet_leaf_119_clk),
    .D(net535),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _13896_ (.CLK(clknet_leaf_120_clk),
    .D(net2149),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _13897_ (.CLK(clknet_leaf_175_clk),
    .D(_00126_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _13898_ (.CLK(clknet_leaf_175_clk),
    .D(_00127_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13899_ (.CLK(clknet_leaf_175_clk),
    .D(_00128_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13900_ (.CLK(clknet_leaf_175_clk),
    .D(_00129_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13901_ (.CLK(clknet_leaf_175_clk),
    .D(_00130_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13902_ (.CLK(clknet_leaf_175_clk),
    .D(_00131_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13903_ (.CLK(clknet_leaf_175_clk),
    .D(_00132_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13904_ (.CLK(clknet_leaf_24_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13905_ (.CLK(clknet_leaf_24_clk),
    .D(net1054),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13906_ (.CLK(clknet_leaf_24_clk),
    .D(net1950),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13907_ (.CLK(clknet_leaf_120_clk),
    .D(net68),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13908_ (.CLK(clknet_leaf_185_clk),
    .D(_00006_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _13909_ (.CLK(clknet_leaf_184_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13910_ (.CLK(clknet_leaf_188_clk),
    .D(net2941),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13911_ (.CLK(clknet_leaf_188_clk),
    .D(net3019),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13912_ (.CLK(clknet_leaf_188_clk),
    .D(net3035),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13913_ (.CLK(clknet_leaf_182_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13914_ (.CLK(clknet_leaf_184_clk),
    .D(net3060),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13915_ (.CLK(clknet_leaf_183_clk),
    .D(net2300),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13916_ (.CLK(clknet_leaf_183_clk),
    .D(net3037),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13917_ (.CLK(clknet_leaf_184_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13918_ (.CLK(clknet_leaf_188_clk),
    .D(net2952),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13919_ (.CLK(clknet_leaf_188_clk),
    .D(net3028),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13920_ (.CLK(clknet_leaf_188_clk),
    .D(net3024),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13921_ (.CLK(clknet_leaf_175_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13922_ (.CLK(clknet_leaf_184_clk),
    .D(net3121),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13923_ (.CLK(clknet_leaf_184_clk),
    .D(net3101),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13924_ (.CLK(clknet_leaf_182_clk),
    .D(net2970),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13925_ (.CLK(clknet_leaf_2_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13926_ (.CLK(clknet_leaf_2_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13927_ (.CLK(clknet_leaf_1_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13928_ (.CLK(clknet_leaf_1_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13929_ (.CLK(clknet_leaf_1_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13930_ (.CLK(clknet_leaf_1_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13931_ (.CLK(clknet_leaf_1_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13932_ (.CLK(clknet_leaf_0_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13933_ (.CLK(clknet_leaf_3_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13934_ (.CLK(clknet_leaf_3_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13935_ (.CLK(clknet_leaf_4_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13936_ (.CLK(clknet_leaf_3_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13937_ (.CLK(clknet_leaf_2_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13938_ (.CLK(clknet_leaf_2_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13939_ (.CLK(clknet_leaf_2_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13940_ (.CLK(clknet_leaf_2_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13941_ (.CLK(clknet_leaf_187_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13942_ (.CLK(clknet_leaf_187_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13943_ (.CLK(clknet_leaf_188_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13944_ (.CLK(clknet_leaf_0_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13945_ (.CLK(clknet_leaf_0_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13946_ (.CLK(clknet_leaf_190_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13947_ (.CLK(clknet_leaf_190_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13948_ (.CLK(clknet_leaf_190_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13949_ (.CLK(clknet_leaf_0_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13950_ (.CLK(clknet_leaf_1_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13951_ (.CLK(clknet_leaf_3_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13952_ (.CLK(clknet_leaf_3_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13953_ (.CLK(clknet_leaf_0_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13954_ (.CLK(clknet_leaf_0_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13955_ (.CLK(clknet_leaf_0_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13956_ (.CLK(clknet_leaf_187_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13957_ (.CLK(clknet_leaf_18_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _13958_ (.CLK(clknet_leaf_5_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _13959_ (.CLK(clknet_leaf_5_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _13960_ (.CLK(clknet_leaf_186_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _13961_ (.CLK(clknet_leaf_186_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _13962_ (.CLK(clknet_leaf_186_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _13963_ (.CLK(clknet_leaf_187_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _13964_ (.CLK(clknet_leaf_187_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _13965_ (.CLK(clknet_leaf_4_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _13966_ (.CLK(clknet_leaf_5_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _13967_ (.CLK(clknet_leaf_5_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _13968_ (.CLK(clknet_leaf_5_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _13969_ (.CLK(clknet_leaf_167_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _13970_ (.CLK(clknet_leaf_167_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _13971_ (.CLK(clknet_leaf_167_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _13972_ (.CLK(clknet_leaf_2_clk),
    .D(net2237),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13973_ (.CLK(clknet_leaf_2_clk),
    .D(net2709),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13974_ (.CLK(clknet_leaf_1_clk),
    .D(net2506),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13975_ (.CLK(clknet_leaf_1_clk),
    .D(net2727),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13976_ (.CLK(clknet_leaf_1_clk),
    .D(net1580),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13977_ (.CLK(clknet_leaf_1_clk),
    .D(net2285),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13978_ (.CLK(clknet_leaf_1_clk),
    .D(net1225),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13979_ (.CLK(clknet_leaf_1_clk),
    .D(net490),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13980_ (.CLK(clknet_leaf_3_clk),
    .D(net1233),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13981_ (.CLK(clknet_leaf_3_clk),
    .D(net2467),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13982_ (.CLK(clknet_leaf_3_clk),
    .D(net236),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13983_ (.CLK(clknet_leaf_3_clk),
    .D(net1719),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13984_ (.CLK(clknet_leaf_2_clk),
    .D(net1151),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13985_ (.CLK(clknet_leaf_2_clk),
    .D(net2731),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13986_ (.CLK(clknet_leaf_2_clk),
    .D(net2679),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13987_ (.CLK(clknet_leaf_2_clk),
    .D(net2669),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13988_ (.CLK(clknet_leaf_187_clk),
    .D(net1605),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13989_ (.CLK(clknet_leaf_187_clk),
    .D(net2425),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13990_ (.CLK(clknet_leaf_187_clk),
    .D(net721),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13991_ (.CLK(clknet_leaf_0_clk),
    .D(net2320),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13992_ (.CLK(clknet_leaf_190_clk),
    .D(net710),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13993_ (.CLK(clknet_leaf_190_clk),
    .D(net1160),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13994_ (.CLK(clknet_leaf_190_clk),
    .D(net1898),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13995_ (.CLK(clknet_leaf_190_clk),
    .D(net2816),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13996_ (.CLK(clknet_leaf_0_clk),
    .D(net2575),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13997_ (.CLK(clknet_leaf_0_clk),
    .D(net632),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13998_ (.CLK(clknet_leaf_4_clk),
    .D(net1064),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13999_ (.CLK(clknet_leaf_3_clk),
    .D(net1889),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14000_ (.CLK(clknet_leaf_0_clk),
    .D(net1583),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14001_ (.CLK(clknet_leaf_0_clk),
    .D(net2364),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14002_ (.CLK(clknet_leaf_0_clk),
    .D(net1587),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14003_ (.CLK(clknet_leaf_187_clk),
    .D(net2082),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14004_ (.CLK(clknet_leaf_173_clk),
    .D(net3108),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14005_ (.CLK(clknet_leaf_5_clk),
    .D(net2589),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14006_ (.CLK(clknet_leaf_5_clk),
    .D(net2792),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14007_ (.CLK(clknet_leaf_186_clk),
    .D(net1145),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14008_ (.CLK(clknet_leaf_186_clk),
    .D(net2353),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14009_ (.CLK(clknet_leaf_186_clk),
    .D(net2331),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14010_ (.CLK(clknet_leaf_187_clk),
    .D(net2670),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14011_ (.CLK(clknet_leaf_187_clk),
    .D(net2417),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14012_ (.CLK(clknet_leaf_4_clk),
    .D(net911),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14013_ (.CLK(clknet_leaf_5_clk),
    .D(net2033),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14014_ (.CLK(clknet_leaf_5_clk),
    .D(net2232),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14015_ (.CLK(clknet_leaf_4_clk),
    .D(net986),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14016_ (.CLK(clknet_leaf_168_clk),
    .D(net114),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14017_ (.CLK(clknet_leaf_120_clk),
    .D(net512),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14018_ (.CLK(clknet_leaf_167_clk),
    .D(net1876),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14019_ (.CLK(clknet_leaf_2_clk),
    .D(net2348),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14020_ (.CLK(clknet_leaf_2_clk),
    .D(net2692),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14021_ (.CLK(clknet_leaf_1_clk),
    .D(net2283),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14022_ (.CLK(clknet_leaf_1_clk),
    .D(net1511),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14023_ (.CLK(clknet_leaf_1_clk),
    .D(net2267),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14024_ (.CLK(clknet_leaf_1_clk),
    .D(net1223),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14025_ (.CLK(clknet_leaf_1_clk),
    .D(net1624),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14026_ (.CLK(clknet_leaf_1_clk),
    .D(net1255),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14027_ (.CLK(clknet_leaf_3_clk),
    .D(net2814),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14028_ (.CLK(clknet_leaf_3_clk),
    .D(net1259),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14029_ (.CLK(clknet_leaf_4_clk),
    .D(net819),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14030_ (.CLK(clknet_leaf_3_clk),
    .D(net1200),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14031_ (.CLK(clknet_leaf_2_clk),
    .D(net1183),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14032_ (.CLK(clknet_leaf_2_clk),
    .D(net2708),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14033_ (.CLK(clknet_leaf_2_clk),
    .D(net1930),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14034_ (.CLK(clknet_leaf_2_clk),
    .D(net1263),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14035_ (.CLK(clknet_leaf_187_clk),
    .D(net1854),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14036_ (.CLK(clknet_leaf_188_clk),
    .D(net732),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14037_ (.CLK(clknet_leaf_188_clk),
    .D(net647),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14038_ (.CLK(clknet_leaf_0_clk),
    .D(net2624),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14039_ (.CLK(clknet_leaf_190_clk),
    .D(net2180),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14040_ (.CLK(clknet_leaf_190_clk),
    .D(net2438),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14041_ (.CLK(clknet_leaf_190_clk),
    .D(net1216),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14042_ (.CLK(clknet_leaf_190_clk),
    .D(net2060),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14043_ (.CLK(clknet_leaf_0_clk),
    .D(net1524),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14044_ (.CLK(clknet_leaf_3_clk),
    .D(net563),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14045_ (.CLK(clknet_leaf_4_clk),
    .D(net1021),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14046_ (.CLK(clknet_leaf_3_clk),
    .D(net2179),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14047_ (.CLK(clknet_leaf_0_clk),
    .D(net1124),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14048_ (.CLK(clknet_leaf_0_clk),
    .D(net2424),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14049_ (.CLK(clknet_leaf_0_clk),
    .D(net2105),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14050_ (.CLK(clknet_leaf_187_clk),
    .D(net1968),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14051_ (.CLK(clknet_leaf_173_clk),
    .D(net1942),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14052_ (.CLK(clknet_leaf_5_clk),
    .D(net2573),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14053_ (.CLK(clknet_leaf_5_clk),
    .D(net2211),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14054_ (.CLK(clknet_leaf_186_clk),
    .D(net2637),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14055_ (.CLK(clknet_leaf_186_clk),
    .D(net1205),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14056_ (.CLK(clknet_leaf_186_clk),
    .D(net1608),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14057_ (.CLK(clknet_leaf_187_clk),
    .D(net2077),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14058_ (.CLK(clknet_leaf_187_clk),
    .D(net2730),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14059_ (.CLK(clknet_leaf_4_clk),
    .D(net1058),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14060_ (.CLK(clknet_leaf_5_clk),
    .D(net1431),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14061_ (.CLK(clknet_leaf_5_clk),
    .D(net1380),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14062_ (.CLK(clknet_leaf_4_clk),
    .D(net1247),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14063_ (.CLK(clknet_leaf_168_clk),
    .D(net2366),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14064_ (.CLK(clknet_leaf_120_clk),
    .D(net2458),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14065_ (.CLK(clknet_leaf_167_clk),
    .D(net1314),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14066_ (.CLK(clknet_leaf_1_clk),
    .D(net472),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14067_ (.CLK(clknet_leaf_1_clk),
    .D(net657),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14068_ (.CLK(clknet_leaf_1_clk),
    .D(net2813),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14069_ (.CLK(clknet_leaf_1_clk),
    .D(net1401),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14070_ (.CLK(clknet_leaf_3_clk),
    .D(net693),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14071_ (.CLK(clknet_leaf_1_clk),
    .D(net2158),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14072_ (.CLK(clknet_leaf_1_clk),
    .D(net1256),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14073_ (.CLK(clknet_leaf_1_clk),
    .D(net2241),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14074_ (.CLK(clknet_leaf_3_clk),
    .D(net2289),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14075_ (.CLK(clknet_leaf_4_clk),
    .D(net2147),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14076_ (.CLK(clknet_leaf_4_clk),
    .D(net1074),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14077_ (.CLK(clknet_leaf_4_clk),
    .D(net853),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14078_ (.CLK(clknet_leaf_2_clk),
    .D(net2667),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14079_ (.CLK(clknet_leaf_2_clk),
    .D(net2847),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14080_ (.CLK(clknet_leaf_3_clk),
    .D(net576),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14081_ (.CLK(clknet_leaf_2_clk),
    .D(net2192),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14082_ (.CLK(clknet_leaf_187_clk),
    .D(net1179),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14083_ (.CLK(clknet_leaf_187_clk),
    .D(net730),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14084_ (.CLK(clknet_leaf_188_clk),
    .D(net1804),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14085_ (.CLK(clknet_leaf_0_clk),
    .D(net2124),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14086_ (.CLK(clknet_leaf_190_clk),
    .D(net954),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14087_ (.CLK(clknet_leaf_190_clk),
    .D(net2823),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14088_ (.CLK(clknet_leaf_190_clk),
    .D(net2056),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14089_ (.CLK(clknet_leaf_190_clk),
    .D(net1468),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14090_ (.CLK(clknet_leaf_4_clk),
    .D(net821),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14091_ (.CLK(clknet_leaf_4_clk),
    .D(net818),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14092_ (.CLK(clknet_leaf_4_clk),
    .D(net849),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14093_ (.CLK(clknet_leaf_4_clk),
    .D(net855),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14094_ (.CLK(clknet_leaf_0_clk),
    .D(net990),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14095_ (.CLK(clknet_leaf_0_clk),
    .D(net1895),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14096_ (.CLK(clknet_leaf_0_clk),
    .D(net1443),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14097_ (.CLK(clknet_leaf_188_clk),
    .D(net494),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14098_ (.CLK(clknet_leaf_174_clk),
    .D(net136),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14099_ (.CLK(clknet_leaf_5_clk),
    .D(net1530),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14100_ (.CLK(clknet_leaf_5_clk),
    .D(net1845),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14101_ (.CLK(clknet_leaf_173_clk),
    .D(net694),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14102_ (.CLK(clknet_leaf_186_clk),
    .D(net2115),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14103_ (.CLK(clknet_leaf_186_clk),
    .D(net1616),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14104_ (.CLK(clknet_leaf_186_clk),
    .D(net88),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14105_ (.CLK(clknet_leaf_186_clk),
    .D(net89),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14106_ (.CLK(clknet_leaf_5_clk),
    .D(net222),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14107_ (.CLK(clknet_leaf_5_clk),
    .D(net1590),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14108_ (.CLK(clknet_leaf_5_clk),
    .D(net1962),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14109_ (.CLK(clknet_leaf_5_clk),
    .D(net221),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14110_ (.CLK(clknet_leaf_167_clk),
    .D(net72),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _14111_ (.CLK(clknet_leaf_120_clk),
    .D(net2716),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _14112_ (.CLK(clknet_leaf_120_clk),
    .D(net477),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_4 _14113_ (.CLK(clknet_leaf_186_clk),
    .D(_00133_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _14114_ (.CLK(clknet_leaf_186_clk),
    .D(_00134_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14115_ (.CLK(clknet_leaf_186_clk),
    .D(_00135_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14116_ (.CLK(clknet_leaf_186_clk),
    .D(_00136_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14117_ (.CLK(clknet_leaf_186_clk),
    .D(_00137_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14118_ (.CLK(clknet_leaf_186_clk),
    .D(_00138_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14119_ (.CLK(clknet_leaf_186_clk),
    .D(_00139_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14120_ (.CLK(clknet_leaf_167_clk),
    .D(_00140_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ));
 sky130_fd_sc_hd__dfxtp_1 _14121_ (.CLK(clknet_leaf_168_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14122_ (.CLK(clknet_leaf_168_clk),
    .D(net2338),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14123_ (.CLK(clknet_leaf_168_clk),
    .D(net1128),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14124_ (.CLK(clknet_leaf_167_clk),
    .D(net77),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14125_ (.CLK(clknet_leaf_187_clk),
    .D(_00007_),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _14126_ (.CLK(clknet_leaf_188_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14127_ (.CLK(clknet_leaf_190_clk),
    .D(net3067),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14128_ (.CLK(clknet_leaf_190_clk),
    .D(net3025),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14129_ (.CLK(clknet_leaf_190_clk),
    .D(net3055),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14130_ (.CLK(clknet_leaf_187_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14131_ (.CLK(clknet_leaf_187_clk),
    .D(net3033),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14132_ (.CLK(clknet_leaf_190_clk),
    .D(net2979),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14133_ (.CLK(clknet_leaf_190_clk),
    .D(net3017),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14134_ (.CLK(clknet_leaf_187_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14135_ (.CLK(clknet_leaf_0_clk),
    .D(net3023),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14136_ (.CLK(clknet_leaf_0_clk),
    .D(net3042),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14137_ (.CLK(clknet_leaf_0_clk),
    .D(net3030),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14138_ (.CLK(clknet_leaf_186_clk),
    .D(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14139_ (.CLK(clknet_leaf_4_clk),
    .D(net3113),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14140_ (.CLK(clknet_leaf_187_clk),
    .D(net2962),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14141_ (.CLK(clknet_leaf_187_clk),
    .D(net3095),
    .Q(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_4 _14142_ (.CLK(clknet_leaf_180_clk),
    .D(net1505),
    .Q(\c.genblk1.genblk1.subs.c0.cfg_i_q[0] ));
 sky130_fd_sc_hd__dfxtp_4 _14143_ (.CLK(clknet_leaf_155_clk),
    .D(net1434),
    .Q(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14144_ (.CLK(clknet_leaf_119_clk),
    .D(net2966),
    .Q(\c.genblk1.genblk1.subs.c0.cfg_i_q[2] ));
 sky130_fd_sc_hd__dfxtp_4 _14145_ (.CLK(clknet_leaf_152_clk),
    .D(net960),
    .Q(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ));
 sky130_fd_sc_hd__dfxtp_4 _14146_ (.CLK(clknet_leaf_146_clk),
    .D(net213),
    .Q(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14147_ (.CLK(clknet_leaf_183_clk),
    .D(net727),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.m[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14148_ (.CLK(clknet_leaf_183_clk),
    .D(net1602),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.m[1] ));
 sky130_fd_sc_hd__dfxtp_4 _14149_ (.CLK(clknet_leaf_189_clk),
    .D(net832),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ));
 sky130_fd_sc_hd__dfxtp_4 _14150_ (.CLK(clknet_leaf_190_clk),
    .D(net1197),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.rst ));
 sky130_fd_sc_hd__dfxtp_1 _14151_ (.CLK(clknet_leaf_8_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14152_ (.CLK(clknet_leaf_3_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14153_ (.CLK(clknet_leaf_2_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14154_ (.CLK(clknet_leaf_3_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14155_ (.CLK(clknet_leaf_8_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14156_ (.CLK(clknet_leaf_7_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14157_ (.CLK(clknet_leaf_9_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14158_ (.CLK(clknet_leaf_8_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14159_ (.CLK(clknet_leaf_20_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14160_ (.CLK(clknet_leaf_18_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14161_ (.CLK(clknet_leaf_172_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14162_ (.CLK(clknet_leaf_173_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14163_ (.CLK(clknet_leaf_8_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14164_ (.CLK(clknet_leaf_2_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14165_ (.CLK(clknet_leaf_8_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14166_ (.CLK(clknet_leaf_8_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14167_ (.CLK(clknet_leaf_18_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14168_ (.CLK(clknet_leaf_18_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14169_ (.CLK(clknet_leaf_172_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14170_ (.CLK(clknet_leaf_173_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14171_ (.CLK(clknet_leaf_6_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14172_ (.CLK(clknet_leaf_6_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14173_ (.CLK(clknet_leaf_4_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14174_ (.CLK(clknet_leaf_7_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14175_ (.CLK(clknet_leaf_19_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14176_ (.CLK(clknet_leaf_18_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14177_ (.CLK(clknet_leaf_172_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14178_ (.CLK(clknet_leaf_173_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14179_ (.CLK(clknet_leaf_7_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14180_ (.CLK(clknet_leaf_7_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14181_ (.CLK(clknet_leaf_7_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14182_ (.CLK(clknet_leaf_6_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14183_ (.CLK(clknet_leaf_19_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14184_ (.CLK(clknet_leaf_22_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14185_ (.CLK(clknet_leaf_22_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14186_ (.CLK(clknet_leaf_22_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14187_ (.CLK(clknet_leaf_172_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14188_ (.CLK(clknet_leaf_169_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14189_ (.CLK(clknet_leaf_22_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14190_ (.CLK(clknet_leaf_22_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14191_ (.CLK(clknet_leaf_19_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14192_ (.CLK(clknet_leaf_19_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14193_ (.CLK(clknet_leaf_172_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14194_ (.CLK(clknet_leaf_172_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14195_ (.CLK(clknet_leaf_23_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14196_ (.CLK(clknet_leaf_23_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14197_ (.CLK(clknet_leaf_23_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14198_ (.CLK(clknet_leaf_8_clk),
    .D(net1931),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14199_ (.CLK(clknet_leaf_7_clk),
    .D(net144),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14200_ (.CLK(clknet_leaf_8_clk),
    .D(net427),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14201_ (.CLK(clknet_leaf_3_clk),
    .D(net2287),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14202_ (.CLK(clknet_leaf_8_clk),
    .D(net2043),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14203_ (.CLK(clknet_leaf_7_clk),
    .D(net2732),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14204_ (.CLK(clknet_leaf_9_clk),
    .D(net2258),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14205_ (.CLK(clknet_leaf_9_clk),
    .D(net125),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14206_ (.CLK(clknet_leaf_19_clk),
    .D(net233),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14207_ (.CLK(clknet_leaf_18_clk),
    .D(net2280),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14208_ (.CLK(clknet_leaf_172_clk),
    .D(net1809),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14209_ (.CLK(clknet_leaf_173_clk),
    .D(net1317),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14210_ (.CLK(clknet_leaf_8_clk),
    .D(net2887),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14211_ (.CLK(clknet_leaf_8_clk),
    .D(net433),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14212_ (.CLK(clknet_leaf_8_clk),
    .D(net2245),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14213_ (.CLK(clknet_leaf_8_clk),
    .D(net1298),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14214_ (.CLK(clknet_leaf_18_clk),
    .D(net1614),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14215_ (.CLK(clknet_leaf_18_clk),
    .D(net2139),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14216_ (.CLK(clknet_leaf_172_clk),
    .D(net1628),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14217_ (.CLK(clknet_leaf_173_clk),
    .D(net1254),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14218_ (.CLK(clknet_leaf_5_clk),
    .D(net607),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14219_ (.CLK(clknet_leaf_7_clk),
    .D(net736),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14220_ (.CLK(clknet_leaf_6_clk),
    .D(net103),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14221_ (.CLK(clknet_leaf_7_clk),
    .D(net1192),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14222_ (.CLK(clknet_leaf_172_clk),
    .D(net505),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14223_ (.CLK(clknet_leaf_18_clk),
    .D(net2206),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14224_ (.CLK(clknet_leaf_172_clk),
    .D(net2805),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14225_ (.CLK(clknet_leaf_173_clk),
    .D(net2705),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14226_ (.CLK(clknet_leaf_7_clk),
    .D(net2207),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14227_ (.CLK(clknet_leaf_7_clk),
    .D(net984),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14228_ (.CLK(clknet_leaf_6_clk),
    .D(net330),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14229_ (.CLK(clknet_leaf_6_clk),
    .D(net2843),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14230_ (.CLK(clknet_leaf_19_clk),
    .D(net2893),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14231_ (.CLK(clknet_leaf_22_clk),
    .D(net2398),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14232_ (.CLK(clknet_leaf_19_clk),
    .D(net643),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14233_ (.CLK(clknet_leaf_22_clk),
    .D(net2446),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14234_ (.CLK(clknet_leaf_169_clk),
    .D(net562),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14235_ (.CLK(clknet_leaf_169_clk),
    .D(net2157),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14236_ (.CLK(clknet_leaf_169_clk),
    .D(net599),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14237_ (.CLK(clknet_leaf_22_clk),
    .D(net1419),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14238_ (.CLK(clknet_leaf_19_clk),
    .D(net2359),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14239_ (.CLK(clknet_leaf_19_clk),
    .D(net2504),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14240_ (.CLK(clknet_leaf_172_clk),
    .D(net2912),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14241_ (.CLK(clknet_leaf_172_clk),
    .D(net2047),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14242_ (.CLK(clknet_leaf_23_clk),
    .D(net1257),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14243_ (.CLK(clknet_leaf_23_clk),
    .D(net1236),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14244_ (.CLK(clknet_leaf_23_clk),
    .D(net2483),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14245_ (.CLK(clknet_leaf_8_clk),
    .D(net2329),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14246_ (.CLK(clknet_leaf_3_clk),
    .D(net366),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14247_ (.CLK(clknet_leaf_3_clk),
    .D(net684),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14248_ (.CLK(clknet_leaf_3_clk),
    .D(net1897),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14249_ (.CLK(clknet_leaf_8_clk),
    .D(net1290),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14250_ (.CLK(clknet_leaf_8_clk),
    .D(net318),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14251_ (.CLK(clknet_leaf_9_clk),
    .D(net1309),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14252_ (.CLK(clknet_leaf_9_clk),
    .D(net1382),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14253_ (.CLK(clknet_leaf_20_clk),
    .D(net792),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14254_ (.CLK(clknet_leaf_18_clk),
    .D(net2789),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14255_ (.CLK(clknet_leaf_172_clk),
    .D(net1353),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14256_ (.CLK(clknet_leaf_173_clk),
    .D(net1637),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14257_ (.CLK(clknet_leaf_8_clk),
    .D(net1746),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14258_ (.CLK(clknet_leaf_2_clk),
    .D(net724),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14259_ (.CLK(clknet_leaf_8_clk),
    .D(net2690),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14260_ (.CLK(clknet_leaf_8_clk),
    .D(net2482),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14261_ (.CLK(clknet_leaf_173_clk),
    .D(net3117),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14262_ (.CLK(clknet_leaf_18_clk),
    .D(net1734),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14263_ (.CLK(clknet_leaf_172_clk),
    .D(net2648),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14264_ (.CLK(clknet_leaf_173_clk),
    .D(net1467),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14265_ (.CLK(clknet_leaf_6_clk),
    .D(net123),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14266_ (.CLK(clknet_leaf_6_clk),
    .D(net285),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14267_ (.CLK(clknet_leaf_6_clk),
    .D(net1111),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14268_ (.CLK(clknet_leaf_6_clk),
    .D(net287),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14269_ (.CLK(clknet_leaf_172_clk),
    .D(net1343),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14270_ (.CLK(clknet_leaf_18_clk),
    .D(net1949),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14271_ (.CLK(clknet_leaf_172_clk),
    .D(net2818),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14272_ (.CLK(clknet_leaf_173_clk),
    .D(net2260),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14273_ (.CLK(clknet_leaf_7_clk),
    .D(net1494),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14274_ (.CLK(clknet_leaf_7_clk),
    .D(net1654),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14275_ (.CLK(clknet_leaf_6_clk),
    .D(net1815),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14276_ (.CLK(clknet_leaf_6_clk),
    .D(net1960),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14277_ (.CLK(clknet_leaf_19_clk),
    .D(net2536),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14278_ (.CLK(clknet_leaf_22_clk),
    .D(net1451),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14279_ (.CLK(clknet_leaf_22_clk),
    .D(net484),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14280_ (.CLK(clknet_leaf_23_clk),
    .D(net523),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14281_ (.CLK(clknet_leaf_172_clk),
    .D(net669),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14282_ (.CLK(clknet_leaf_169_clk),
    .D(net1286),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14283_ (.CLK(clknet_leaf_169_clk),
    .D(net2270),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14284_ (.CLK(clknet_leaf_169_clk),
    .D(net475),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14285_ (.CLK(clknet_leaf_19_clk),
    .D(net1313),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14286_ (.CLK(clknet_leaf_19_clk),
    .D(net2510),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14287_ (.CLK(clknet_leaf_171_clk),
    .D(net501),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14288_ (.CLK(clknet_leaf_172_clk),
    .D(net2341),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14289_ (.CLK(clknet_leaf_168_clk),
    .D(net581),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14290_ (.CLK(clknet_leaf_23_clk),
    .D(net1342),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14291_ (.CLK(clknet_leaf_23_clk),
    .D(net2177),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14292_ (.CLK(clknet_leaf_8_clk),
    .D(net2090),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14293_ (.CLK(clknet_leaf_7_clk),
    .D(net146),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14294_ (.CLK(clknet_leaf_8_clk),
    .D(net555),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14295_ (.CLK(clknet_leaf_3_clk),
    .D(net2014),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14296_ (.CLK(clknet_leaf_8_clk),
    .D(net2256),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14297_ (.CLK(clknet_leaf_7_clk),
    .D(net143),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14298_ (.CLK(clknet_leaf_9_clk),
    .D(net1378),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14299_ (.CLK(clknet_leaf_9_clk),
    .D(net2150),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14300_ (.CLK(clknet_leaf_19_clk),
    .D(net269),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14301_ (.CLK(clknet_leaf_18_clk),
    .D(net2892),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14302_ (.CLK(clknet_leaf_171_clk),
    .D(net766),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14303_ (.CLK(clknet_leaf_172_clk),
    .D(net546),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14304_ (.CLK(clknet_leaf_8_clk),
    .D(net1445),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14305_ (.CLK(clknet_leaf_2_clk),
    .D(net1159),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14306_ (.CLK(clknet_leaf_8_clk),
    .D(net2492),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14307_ (.CLK(clknet_leaf_8_clk),
    .D(net2910),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14308_ (.CLK(clknet_leaf_18_clk),
    .D(net41),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14309_ (.CLK(clknet_leaf_173_clk),
    .D(net3114),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14310_ (.CLK(clknet_leaf_172_clk),
    .D(net1666),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14311_ (.CLK(clknet_leaf_172_clk),
    .D(net479),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14312_ (.CLK(clknet_leaf_6_clk),
    .D(net1076),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14313_ (.CLK(clknet_leaf_6_clk),
    .D(net1084),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14314_ (.CLK(clknet_leaf_6_clk),
    .D(net1376),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14315_ (.CLK(clknet_leaf_6_clk),
    .D(net1751),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14316_ (.CLK(clknet_leaf_172_clk),
    .D(net1836),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14317_ (.CLK(clknet_leaf_18_clk),
    .D(net2205),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14318_ (.CLK(clknet_leaf_171_clk),
    .D(net725),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14319_ (.CLK(clknet_leaf_173_clk),
    .D(net2831),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14320_ (.CLK(clknet_leaf_6_clk),
    .D(net268),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14321_ (.CLK(clknet_leaf_7_clk),
    .D(net2900),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14322_ (.CLK(clknet_leaf_6_clk),
    .D(net2153),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14323_ (.CLK(clknet_leaf_6_clk),
    .D(net1227),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14324_ (.CLK(clknet_leaf_19_clk),
    .D(net2324),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14325_ (.CLK(clknet_leaf_169_clk),
    .D(net630),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14326_ (.CLK(clknet_leaf_22_clk),
    .D(net2096),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14327_ (.CLK(clknet_leaf_169_clk),
    .D(net548),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14328_ (.CLK(clknet_leaf_169_clk),
    .D(net570),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14329_ (.CLK(clknet_leaf_169_clk),
    .D(net2128),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14330_ (.CLK(clknet_leaf_169_clk),
    .D(net2456),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14331_ (.CLK(clknet_leaf_169_clk),
    .D(net2556),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14332_ (.CLK(clknet_leaf_19_clk),
    .D(net1828),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14333_ (.CLK(clknet_leaf_19_clk),
    .D(net2600),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14334_ (.CLK(clknet_leaf_172_clk),
    .D(net706),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14335_ (.CLK(clknet_leaf_172_clk),
    .D(net2361),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14336_ (.CLK(clknet_leaf_168_clk),
    .D(net2457),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _14337_ (.CLK(clknet_leaf_23_clk),
    .D(net1476),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _14338_ (.CLK(clknet_leaf_23_clk),
    .D(net1607),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _14339_ (.CLK(clknet_leaf_20_clk),
    .D(_00141_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _14340_ (.CLK(clknet_leaf_18_clk),
    .D(net3183),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14341_ (.CLK(clknet_leaf_17_clk),
    .D(_00143_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14342_ (.CLK(clknet_leaf_17_clk),
    .D(_00144_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14343_ (.CLK(clknet_leaf_18_clk),
    .D(net3671),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14344_ (.CLK(clknet_leaf_19_clk),
    .D(_00146_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14345_ (.CLK(clknet_leaf_19_clk),
    .D(_00147_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14346_ (.CLK(clknet_leaf_63_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14347_ (.CLK(clknet_leaf_67_clk),
    .D(net471),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14348_ (.CLK(clknet_leaf_67_clk),
    .D(net2395),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14349_ (.CLK(clknet_leaf_67_clk),
    .D(net1766),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14350_ (.CLK(clknet_leaf_6_clk),
    .D(_00000_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _14351_ (.CLK(clknet_leaf_18_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14352_ (.CLK(clknet_leaf_17_clk),
    .D(net3165),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14353_ (.CLK(clknet_leaf_17_clk),
    .D(net3086),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14354_ (.CLK(clknet_leaf_18_clk),
    .D(net113),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14355_ (.CLK(clknet_leaf_18_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14356_ (.CLK(clknet_leaf_18_clk),
    .D(net3029),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14357_ (.CLK(clknet_leaf_18_clk),
    .D(net3027),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14358_ (.CLK(clknet_leaf_5_clk),
    .D(net3178),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14359_ (.CLK(clknet_leaf_17_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14360_ (.CLK(clknet_leaf_5_clk),
    .D(net3001),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14361_ (.CLK(clknet_leaf_5_clk),
    .D(net3034),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14362_ (.CLK(clknet_leaf_5_clk),
    .D(net3058),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14363_ (.CLK(clknet_leaf_18_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14364_ (.CLK(clknet_leaf_6_clk),
    .D(net3220),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14365_ (.CLK(clknet_leaf_5_clk),
    .D(net3053),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14366_ (.CLK(clknet_leaf_18_clk),
    .D(net66),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14367_ (.CLK(clknet_leaf_11_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14368_ (.CLK(clknet_leaf_11_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14369_ (.CLK(clknet_leaf_10_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14370_ (.CLK(clknet_leaf_11_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14371_ (.CLK(clknet_leaf_11_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14372_ (.CLK(clknet_leaf_11_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14373_ (.CLK(clknet_leaf_11_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14374_ (.CLK(clknet_leaf_12_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14375_ (.CLK(clknet_leaf_15_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14376_ (.CLK(clknet_leaf_14_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14377_ (.CLK(clknet_leaf_14_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14378_ (.CLK(clknet_leaf_14_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14379_ (.CLK(clknet_leaf_14_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14380_ (.CLK(clknet_leaf_10_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14381_ (.CLK(clknet_leaf_13_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14382_ (.CLK(clknet_leaf_13_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14383_ (.CLK(clknet_leaf_17_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14384_ (.CLK(clknet_leaf_17_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14385_ (.CLK(clknet_leaf_16_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14386_ (.CLK(clknet_leaf_16_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14387_ (.CLK(clknet_leaf_9_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14388_ (.CLK(clknet_leaf_9_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14389_ (.CLK(clknet_leaf_9_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14390_ (.CLK(clknet_leaf_9_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14391_ (.CLK(clknet_leaf_17_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14392_ (.CLK(clknet_leaf_10_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14393_ (.CLK(clknet_leaf_13_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14394_ (.CLK(clknet_leaf_16_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14395_ (.CLK(clknet_leaf_10_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14396_ (.CLK(clknet_leaf_9_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14397_ (.CLK(clknet_leaf_9_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14398_ (.CLK(clknet_leaf_9_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14399_ (.CLK(clknet_leaf_21_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14400_ (.CLK(clknet_leaf_19_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14401_ (.CLK(clknet_leaf_22_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14402_ (.CLK(clknet_leaf_21_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14403_ (.CLK(clknet_leaf_22_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14404_ (.CLK(clknet_leaf_23_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14405_ (.CLK(clknet_leaf_20_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14406_ (.CLK(clknet_leaf_19_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14407_ (.CLK(clknet_leaf_20_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14408_ (.CLK(clknet_leaf_20_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14409_ (.CLK(clknet_leaf_15_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14410_ (.CLK(clknet_leaf_15_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14411_ (.CLK(clknet_leaf_23_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14412_ (.CLK(clknet_leaf_23_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14413_ (.CLK(clknet_leaf_24_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14414_ (.CLK(clknet_leaf_11_clk),
    .D(net2820),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14415_ (.CLK(clknet_leaf_11_clk),
    .D(net1118),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14416_ (.CLK(clknet_leaf_11_clk),
    .D(net770),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14417_ (.CLK(clknet_leaf_11_clk),
    .D(net2091),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14418_ (.CLK(clknet_leaf_12_clk),
    .D(net692),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14419_ (.CLK(clknet_leaf_11_clk),
    .D(net2185),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14420_ (.CLK(clknet_leaf_11_clk),
    .D(net1659),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14421_ (.CLK(clknet_leaf_12_clk),
    .D(net1191),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14422_ (.CLK(clknet_leaf_15_clk),
    .D(net2461),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14423_ (.CLK(clknet_leaf_16_clk),
    .D(net889),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14424_ (.CLK(clknet_leaf_14_clk),
    .D(net2653),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14425_ (.CLK(clknet_leaf_13_clk),
    .D(net493),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14426_ (.CLK(clknet_leaf_13_clk),
    .D(net644),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14427_ (.CLK(clknet_leaf_10_clk),
    .D(net2517),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14428_ (.CLK(clknet_leaf_13_clk),
    .D(net2945),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14429_ (.CLK(clknet_leaf_13_clk),
    .D(net2923),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14430_ (.CLK(clknet_leaf_17_clk),
    .D(net2269),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14431_ (.CLK(clknet_leaf_17_clk),
    .D(net2689),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14432_ (.CLK(clknet_leaf_17_clk),
    .D(net191),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14433_ (.CLK(clknet_leaf_16_clk),
    .D(net924),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14434_ (.CLK(clknet_leaf_10_clk),
    .D(net461),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14435_ (.CLK(clknet_leaf_9_clk),
    .D(net1733),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14436_ (.CLK(clknet_leaf_11_clk),
    .D(net642),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14437_ (.CLK(clknet_leaf_9_clk),
    .D(net2259),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14438_ (.CLK(clknet_leaf_17_clk),
    .D(net2365),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14439_ (.CLK(clknet_leaf_13_clk),
    .D(net726),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14440_ (.CLK(clknet_leaf_16_clk),
    .D(net2203),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14441_ (.CLK(clknet_leaf_16_clk),
    .D(net1330),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14442_ (.CLK(clknet_leaf_10_clk),
    .D(net1508),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14443_ (.CLK(clknet_leaf_10_clk),
    .D(net385),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14444_ (.CLK(clknet_leaf_9_clk),
    .D(net2265),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14445_ (.CLK(clknet_leaf_9_clk),
    .D(net2295),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14446_ (.CLK(clknet_leaf_21_clk),
    .D(net2336),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14447_ (.CLK(clknet_leaf_19_clk),
    .D(net2799),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14448_ (.CLK(clknet_leaf_22_clk),
    .D(net1945),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14449_ (.CLK(clknet_leaf_22_clk),
    .D(net280),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14450_ (.CLK(clknet_leaf_22_clk),
    .D(net1454),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14451_ (.CLK(clknet_leaf_22_clk),
    .D(net656),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14452_ (.CLK(clknet_leaf_21_clk),
    .D(net337),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14453_ (.CLK(clknet_leaf_19_clk),
    .D(net2344),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14454_ (.CLK(clknet_leaf_20_clk),
    .D(net982),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14455_ (.CLK(clknet_leaf_20_clk),
    .D(net962),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14456_ (.CLK(clknet_leaf_15_clk),
    .D(net1155),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14457_ (.CLK(clknet_leaf_15_clk),
    .D(net1135),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14458_ (.CLK(clknet_leaf_23_clk),
    .D(net2000),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14459_ (.CLK(clknet_leaf_23_clk),
    .D(net1597),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14460_ (.CLK(clknet_leaf_24_clk),
    .D(net1046),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14461_ (.CLK(clknet_leaf_11_clk),
    .D(net2222),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14462_ (.CLK(clknet_leaf_11_clk),
    .D(net1146),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14463_ (.CLK(clknet_leaf_10_clk),
    .D(net322),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14464_ (.CLK(clknet_leaf_11_clk),
    .D(net2688),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14465_ (.CLK(clknet_leaf_11_clk),
    .D(net344),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14466_ (.CLK(clknet_leaf_11_clk),
    .D(net2089),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14467_ (.CLK(clknet_leaf_11_clk),
    .D(net2521),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14468_ (.CLK(clknet_leaf_12_clk),
    .D(net2092),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14469_ (.CLK(clknet_leaf_15_clk),
    .D(net2172),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14470_ (.CLK(clknet_leaf_16_clk),
    .D(net856),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14471_ (.CLK(clknet_leaf_14_clk),
    .D(net2473),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14472_ (.CLK(clknet_leaf_14_clk),
    .D(net515),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14473_ (.CLK(clknet_leaf_14_clk),
    .D(net467),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14474_ (.CLK(clknet_leaf_10_clk),
    .D(net1625),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14475_ (.CLK(clknet_leaf_13_clk),
    .D(net1754),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14476_ (.CLK(clknet_leaf_13_clk),
    .D(net1752),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14477_ (.CLK(clknet_leaf_17_clk),
    .D(net2038),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14478_ (.CLK(clknet_leaf_17_clk),
    .D(net1646),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14479_ (.CLK(clknet_leaf_17_clk),
    .D(net1921),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14480_ (.CLK(clknet_leaf_17_clk),
    .D(net202),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14481_ (.CLK(clknet_leaf_10_clk),
    .D(net2850),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14482_ (.CLK(clknet_leaf_9_clk),
    .D(net1316),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14483_ (.CLK(clknet_leaf_11_clk),
    .D(net1562),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14484_ (.CLK(clknet_leaf_9_clk),
    .D(net2340),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14485_ (.CLK(clknet_leaf_17_clk),
    .D(net2240),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14486_ (.CLK(clknet_leaf_13_clk),
    .D(net1642),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14487_ (.CLK(clknet_leaf_13_clk),
    .D(net184),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14488_ (.CLK(clknet_leaf_16_clk),
    .D(net920),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14489_ (.CLK(clknet_leaf_7_clk),
    .D(net778),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14490_ (.CLK(clknet_leaf_10_clk),
    .D(net2770),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14491_ (.CLK(clknet_leaf_9_clk),
    .D(net2176),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14492_ (.CLK(clknet_leaf_9_clk),
    .D(net1868),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14493_ (.CLK(clknet_leaf_21_clk),
    .D(net1001),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14494_ (.CLK(clknet_leaf_19_clk),
    .D(net2160),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14495_ (.CLK(clknet_leaf_22_clk),
    .D(net2286),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14496_ (.CLK(clknet_leaf_22_clk),
    .D(net2567),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14497_ (.CLK(clknet_leaf_23_clk),
    .D(net603),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14498_ (.CLK(clknet_leaf_22_clk),
    .D(net1555),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14499_ (.CLK(clknet_leaf_20_clk),
    .D(net734),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14500_ (.CLK(clknet_leaf_19_clk),
    .D(net1905),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14501_ (.CLK(clknet_leaf_20_clk),
    .D(net980),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14502_ (.CLK(clknet_leaf_20_clk),
    .D(net2214),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14503_ (.CLK(clknet_leaf_15_clk),
    .D(net1169),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14504_ (.CLK(clknet_leaf_20_clk),
    .D(net283),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14505_ (.CLK(clknet_leaf_23_clk),
    .D(net1279),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14506_ (.CLK(clknet_leaf_23_clk),
    .D(net1744),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14507_ (.CLK(clknet_leaf_24_clk),
    .D(net2182),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14508_ (.CLK(clknet_leaf_11_clk),
    .D(net1215),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14509_ (.CLK(clknet_leaf_10_clk),
    .D(net340),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14510_ (.CLK(clknet_leaf_10_clk),
    .D(net1913),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14511_ (.CLK(clknet_leaf_10_clk),
    .D(net375),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14512_ (.CLK(clknet_leaf_11_clk),
    .D(net1117),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14513_ (.CLK(clknet_leaf_11_clk),
    .D(net2112),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14514_ (.CLK(clknet_leaf_11_clk),
    .D(net2711),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14515_ (.CLK(clknet_leaf_13_clk),
    .D(net310),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14516_ (.CLK(clknet_leaf_15_clk),
    .D(net2362),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14517_ (.CLK(clknet_leaf_16_clk),
    .D(net888),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14518_ (.CLK(clknet_leaf_14_clk),
    .D(net1994),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14519_ (.CLK(clknet_leaf_14_clk),
    .D(net1544),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14520_ (.CLK(clknet_leaf_14_clk),
    .D(net1834),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14521_ (.CLK(clknet_leaf_13_clk),
    .D(net686),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14522_ (.CLK(clknet_leaf_13_clk),
    .D(net1331),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14523_ (.CLK(clknet_leaf_13_clk),
    .D(net1326),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14524_ (.CLK(clknet_leaf_17_clk),
    .D(net1727),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14525_ (.CLK(clknet_leaf_17_clk),
    .D(net2890),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14526_ (.CLK(clknet_leaf_17_clk),
    .D(net2162),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14527_ (.CLK(clknet_leaf_16_clk),
    .D(net1584),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14528_ (.CLK(clknet_leaf_10_clk),
    .D(net1546),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14529_ (.CLK(clknet_leaf_10_clk),
    .D(net440),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14530_ (.CLK(clknet_leaf_10_clk),
    .D(net365),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14531_ (.CLK(clknet_leaf_9_clk),
    .D(net2371),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14532_ (.CLK(clknet_leaf_17_clk),
    .D(net1057),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14533_ (.CLK(clknet_leaf_13_clk),
    .D(net2367),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14534_ (.CLK(clknet_leaf_13_clk),
    .D(net1444),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14535_ (.CLK(clknet_leaf_16_clk),
    .D(net1615),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14536_ (.CLK(clknet_leaf_7_clk),
    .D(net991),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14537_ (.CLK(clknet_leaf_10_clk),
    .D(net2159),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14538_ (.CLK(clknet_leaf_9_clk),
    .D(net1826),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14539_ (.CLK(clknet_leaf_9_clk),
    .D(net2084),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14540_ (.CLK(clknet_leaf_22_clk),
    .D(net277),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14541_ (.CLK(clknet_leaf_22_clk),
    .D(net491),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14542_ (.CLK(clknet_leaf_23_clk),
    .D(net645),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14543_ (.CLK(clknet_leaf_22_clk),
    .D(net2677),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14544_ (.CLK(clknet_leaf_23_clk),
    .D(net1579),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14545_ (.CLK(clknet_leaf_23_clk),
    .D(net606),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14546_ (.CLK(clknet_leaf_21_clk),
    .D(net326),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14547_ (.CLK(clknet_leaf_19_clk),
    .D(net2076),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14548_ (.CLK(clknet_leaf_20_clk),
    .D(net1341),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14549_ (.CLK(clknet_leaf_20_clk),
    .D(net1012),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14550_ (.CLK(clknet_leaf_15_clk),
    .D(net1297),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14551_ (.CLK(clknet_leaf_20_clk),
    .D(net1358),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14552_ (.CLK(clknet_leaf_24_clk),
    .D(net147),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _14553_ (.CLK(clknet_leaf_24_clk),
    .D(net151),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _14554_ (.CLK(clknet_leaf_24_clk),
    .D(net2252),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _14555_ (.CLK(clknet_leaf_20_clk),
    .D(_00148_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _14556_ (.CLK(clknet_leaf_20_clk),
    .D(_00149_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14557_ (.CLK(clknet_leaf_20_clk),
    .D(_00150_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14558_ (.CLK(clknet_leaf_20_clk),
    .D(_00151_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14559_ (.CLK(clknet_leaf_15_clk),
    .D(_00152_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14560_ (.CLK(clknet_leaf_16_clk),
    .D(_00153_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14561_ (.CLK(clknet_leaf_16_clk),
    .D(_00154_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14562_ (.CLK(clknet_leaf_63_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14563_ (.CLK(clknet_leaf_67_clk),
    .D(net511),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14564_ (.CLK(clknet_leaf_68_clk),
    .D(net521),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14565_ (.CLK(clknet_leaf_68_clk),
    .D(net1969),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14566_ (.CLK(clknet_leaf_17_clk),
    .D(_00001_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _14567_ (.CLK(clknet_leaf_6_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14568_ (.CLK(clknet_leaf_7_clk),
    .D(net2982),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14569_ (.CLK(clknet_leaf_7_clk),
    .D(net3009),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14570_ (.CLK(clknet_leaf_7_clk),
    .D(net3031),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14571_ (.CLK(clknet_leaf_13_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14572_ (.CLK(clknet_leaf_10_clk),
    .D(net2963),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14573_ (.CLK(clknet_leaf_10_clk),
    .D(net3015),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14574_ (.CLK(clknet_leaf_10_clk),
    .D(net3048),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14575_ (.CLK(clknet_leaf_13_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14576_ (.CLK(clknet_leaf_10_clk),
    .D(net2990),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14577_ (.CLK(clknet_leaf_10_clk),
    .D(net3069),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14578_ (.CLK(clknet_leaf_10_clk),
    .D(net3094),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14579_ (.CLK(clknet_leaf_16_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14580_ (.CLK(clknet_leaf_17_clk),
    .D(net2955),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14581_ (.CLK(clknet_leaf_6_clk),
    .D(net3012),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14582_ (.CLK(clknet_leaf_17_clk),
    .D(net2988),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14583_ (.CLK(clknet_leaf_12_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14584_ (.CLK(clknet_leaf_11_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14585_ (.CLK(clknet_leaf_12_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14586_ (.CLK(clknet_leaf_12_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14587_ (.CLK(clknet_leaf_37_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14588_ (.CLK(clknet_leaf_36_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14589_ (.CLK(clknet_leaf_36_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14590_ (.CLK(clknet_leaf_37_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14591_ (.CLK(clknet_leaf_21_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14592_ (.CLK(clknet_leaf_15_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14593_ (.CLK(clknet_leaf_33_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14594_ (.CLK(clknet_leaf_15_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14595_ (.CLK(clknet_leaf_12_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14596_ (.CLK(clknet_leaf_36_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14597_ (.CLK(clknet_leaf_36_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14598_ (.CLK(clknet_leaf_36_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14599_ (.CLK(clknet_leaf_14_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14600_ (.CLK(clknet_leaf_14_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14601_ (.CLK(clknet_leaf_21_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14602_ (.CLK(clknet_leaf_15_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14603_ (.CLK(clknet_leaf_35_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14604_ (.CLK(clknet_leaf_12_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14605_ (.CLK(clknet_leaf_13_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14606_ (.CLK(clknet_leaf_13_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14607_ (.CLK(clknet_leaf_33_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14608_ (.CLK(clknet_leaf_14_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14609_ (.CLK(clknet_leaf_26_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14610_ (.CLK(clknet_leaf_33_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14611_ (.CLK(clknet_leaf_35_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14612_ (.CLK(clknet_leaf_35_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14613_ (.CLK(clknet_leaf_35_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14614_ (.CLK(clknet_leaf_35_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14615_ (.CLK(clknet_leaf_25_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14616_ (.CLK(clknet_leaf_27_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14617_ (.CLK(clknet_leaf_26_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14618_ (.CLK(clknet_leaf_25_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14619_ (.CLK(clknet_leaf_25_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14620_ (.CLK(clknet_leaf_25_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14621_ (.CLK(clknet_leaf_22_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14622_ (.CLK(clknet_leaf_26_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14623_ (.CLK(clknet_leaf_26_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14624_ (.CLK(clknet_leaf_21_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14625_ (.CLK(clknet_leaf_21_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14626_ (.CLK(clknet_leaf_26_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14627_ (.CLK(clknet_leaf_24_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14628_ (.CLK(clknet_leaf_24_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14629_ (.CLK(clknet_leaf_24_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14630_ (.CLK(clknet_leaf_12_clk),
    .D(net1961),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14631_ (.CLK(clknet_leaf_12_clk),
    .D(net709),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14632_ (.CLK(clknet_leaf_12_clk),
    .D(net1670),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14633_ (.CLK(clknet_leaf_12_clk),
    .D(net1406),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14634_ (.CLK(clknet_leaf_36_clk),
    .D(net587),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14635_ (.CLK(clknet_leaf_36_clk),
    .D(net2668),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14636_ (.CLK(clknet_leaf_36_clk),
    .D(net1686),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14637_ (.CLK(clknet_leaf_36_clk),
    .D(net492),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14638_ (.CLK(clknet_leaf_21_clk),
    .D(net1139),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14639_ (.CLK(clknet_leaf_15_clk),
    .D(net1158),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14640_ (.CLK(clknet_leaf_33_clk),
    .D(net2647),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14641_ (.CLK(clknet_leaf_15_clk),
    .D(net1137),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14642_ (.CLK(clknet_leaf_36_clk),
    .D(net118),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14643_ (.CLK(clknet_leaf_36_clk),
    .D(net2373),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14644_ (.CLK(clknet_leaf_36_clk),
    .D(net1594),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14645_ (.CLK(clknet_leaf_36_clk),
    .D(net2194),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14646_ (.CLK(clknet_leaf_14_clk),
    .D(net1455),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14647_ (.CLK(clknet_leaf_14_clk),
    .D(net2564),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14648_ (.CLK(clknet_leaf_15_clk),
    .D(net106),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14649_ (.CLK(clknet_leaf_15_clk),
    .D(net2542),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14650_ (.CLK(clknet_leaf_36_clk),
    .D(net347),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14651_ (.CLK(clknet_leaf_35_clk),
    .D(net129),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14652_ (.CLK(clknet_leaf_13_clk),
    .D(net2144),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14653_ (.CLK(clknet_leaf_12_clk),
    .D(net707),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14654_ (.CLK(clknet_leaf_33_clk),
    .D(net2577),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14655_ (.CLK(clknet_leaf_15_clk),
    .D(net480),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14656_ (.CLK(clknet_leaf_26_clk),
    .D(net1629),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14657_ (.CLK(clknet_leaf_33_clk),
    .D(net1603),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14658_ (.CLK(clknet_leaf_34_clk),
    .D(net764),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14659_ (.CLK(clknet_leaf_35_clk),
    .D(net1658),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14660_ (.CLK(clknet_leaf_36_clk),
    .D(net352),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14661_ (.CLK(clknet_leaf_35_clk),
    .D(net1979),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14662_ (.CLK(clknet_leaf_25_clk),
    .D(net1997),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14663_ (.CLK(clknet_leaf_28_clk),
    .D(net208),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14664_ (.CLK(clknet_leaf_25_clk),
    .D(net235),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14665_ (.CLK(clknet_leaf_26_clk),
    .D(net846),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14666_ (.CLK(clknet_leaf_25_clk),
    .D(net2030),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14667_ (.CLK(clknet_leaf_25_clk),
    .D(net1785),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14668_ (.CLK(clknet_leaf_23_clk),
    .D(net598),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14669_ (.CLK(clknet_leaf_25_clk),
    .D(net228),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14670_ (.CLK(clknet_leaf_26_clk),
    .D(net971),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14671_ (.CLK(clknet_leaf_21_clk),
    .D(net2781),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14672_ (.CLK(clknet_leaf_21_clk),
    .D(net1047),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14673_ (.CLK(clknet_leaf_26_clk),
    .D(net897),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14674_ (.CLK(clknet_leaf_24_clk),
    .D(net1162),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14675_ (.CLK(clknet_leaf_24_clk),
    .D(net1071),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14676_ (.CLK(clknet_leaf_24_clk),
    .D(net2754),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14677_ (.CLK(clknet_leaf_12_clk),
    .D(net1037),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14678_ (.CLK(clknet_leaf_12_clk),
    .D(net1040),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14679_ (.CLK(clknet_leaf_12_clk),
    .D(net2169),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14680_ (.CLK(clknet_leaf_12_clk),
    .D(net2100),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14681_ (.CLK(clknet_leaf_37_clk),
    .D(net509),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14682_ (.CLK(clknet_leaf_37_clk),
    .D(net464),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14683_ (.CLK(clknet_leaf_36_clk),
    .D(net2197),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14684_ (.CLK(clknet_leaf_37_clk),
    .D(net624),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14685_ (.CLK(clknet_leaf_21_clk),
    .D(net1553),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14686_ (.CLK(clknet_leaf_15_clk),
    .D(net2646),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14687_ (.CLK(clknet_leaf_33_clk),
    .D(net2057),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14688_ (.CLK(clknet_leaf_21_clk),
    .D(net252),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14689_ (.CLK(clknet_leaf_36_clk),
    .D(net2753),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14690_ (.CLK(clknet_leaf_36_clk),
    .D(net1999),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14691_ (.CLK(clknet_leaf_36_clk),
    .D(net2601),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14692_ (.CLK(clknet_leaf_36_clk),
    .D(net1683),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14693_ (.CLK(clknet_leaf_14_clk),
    .D(net2785),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14694_ (.CLK(clknet_leaf_14_clk),
    .D(net2864),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14695_ (.CLK(clknet_leaf_21_clk),
    .D(net250),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14696_ (.CLK(clknet_leaf_15_clk),
    .D(net2067),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14697_ (.CLK(clknet_leaf_12_clk),
    .D(net135),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14698_ (.CLK(clknet_leaf_35_clk),
    .D(net1034),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14699_ (.CLK(clknet_leaf_14_clk),
    .D(net667),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14700_ (.CLK(clknet_leaf_13_clk),
    .D(net303),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14701_ (.CLK(clknet_leaf_33_clk),
    .D(net1481),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14702_ (.CLK(clknet_leaf_15_clk),
    .D(net2744),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14703_ (.CLK(clknet_leaf_26_clk),
    .D(net1007),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14704_ (.CLK(clknet_leaf_33_clk),
    .D(net2277),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14705_ (.CLK(clknet_leaf_34_clk),
    .D(net931),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14706_ (.CLK(clknet_leaf_35_clk),
    .D(net1585),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14707_ (.CLK(clknet_leaf_35_clk),
    .D(net723),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14708_ (.CLK(clknet_leaf_35_clk),
    .D(net2582),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14709_ (.CLK(clknet_leaf_25_clk),
    .D(net1529),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14710_ (.CLK(clknet_leaf_26_clk),
    .D(net812),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14711_ (.CLK(clknet_leaf_26_clk),
    .D(net859),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14712_ (.CLK(clknet_leaf_26_clk),
    .D(net1251),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14713_ (.CLK(clknet_leaf_25_clk),
    .D(net1523),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14714_ (.CLK(clknet_leaf_67_clk),
    .D(net508),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14715_ (.CLK(clknet_leaf_23_clk),
    .D(net1721),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14716_ (.CLK(clknet_leaf_24_clk),
    .D(net695),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14717_ (.CLK(clknet_leaf_26_clk),
    .D(net948),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14718_ (.CLK(clknet_leaf_21_clk),
    .D(net2773),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14719_ (.CLK(clknet_leaf_21_clk),
    .D(net959),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14720_ (.CLK(clknet_leaf_26_clk),
    .D(net2363),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14721_ (.CLK(clknet_leaf_24_clk),
    .D(net1599),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14722_ (.CLK(clknet_leaf_24_clk),
    .D(net2239),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14723_ (.CLK(clknet_leaf_24_clk),
    .D(net1832),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14724_ (.CLK(clknet_leaf_12_clk),
    .D(net2035),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14725_ (.CLK(clknet_leaf_12_clk),
    .D(net1712),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14726_ (.CLK(clknet_leaf_12_clk),
    .D(net1878),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14727_ (.CLK(clknet_leaf_12_clk),
    .D(net1682),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14728_ (.CLK(clknet_leaf_37_clk),
    .D(net2587),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14729_ (.CLK(clknet_leaf_37_clk),
    .D(net2095),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14730_ (.CLK(clknet_leaf_36_clk),
    .D(net1954),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14731_ (.CLK(clknet_leaf_35_clk),
    .D(net601),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14732_ (.CLK(clknet_leaf_21_clk),
    .D(net1413),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14733_ (.CLK(clknet_leaf_15_clk),
    .D(net2138),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14734_ (.CLK(clknet_leaf_33_clk),
    .D(net2154),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14735_ (.CLK(clknet_leaf_21_clk),
    .D(net2026),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14736_ (.CLK(clknet_leaf_36_clk),
    .D(net1940),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14737_ (.CLK(clknet_leaf_36_clk),
    .D(net2439),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14738_ (.CLK(clknet_leaf_36_clk),
    .D(net2930),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14739_ (.CLK(clknet_leaf_36_clk),
    .D(net1327),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14740_ (.CLK(clknet_leaf_14_clk),
    .D(net1373),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14741_ (.CLK(clknet_leaf_14_clk),
    .D(net2616),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14742_ (.CLK(clknet_leaf_21_clk),
    .D(net1193),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14743_ (.CLK(clknet_leaf_15_clk),
    .D(net2188),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14744_ (.CLK(clknet_leaf_35_clk),
    .D(net115),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14745_ (.CLK(clknet_leaf_35_clk),
    .D(net1517),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14746_ (.CLK(clknet_leaf_14_clk),
    .D(net2477),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14747_ (.CLK(clknet_leaf_13_clk),
    .D(net1975),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14748_ (.CLK(clknet_leaf_33_clk),
    .D(net1105),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14749_ (.CLK(clknet_leaf_33_clk),
    .D(net124),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14750_ (.CLK(clknet_leaf_26_clk),
    .D(net1470),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14751_ (.CLK(clknet_leaf_33_clk),
    .D(net1708),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14752_ (.CLK(clknet_leaf_34_clk),
    .D(net1207),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14753_ (.CLK(clknet_leaf_35_clk),
    .D(net1477),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14754_ (.CLK(clknet_leaf_35_clk),
    .D(net1092),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14755_ (.CLK(clknet_leaf_35_clk),
    .D(net2199),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14756_ (.CLK(clknet_leaf_25_clk),
    .D(net2485),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14757_ (.CLK(clknet_leaf_25_clk),
    .D(net227),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14758_ (.CLK(clknet_leaf_26_clk),
    .D(net2009),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14759_ (.CLK(clknet_leaf_25_clk),
    .D(net240),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14760_ (.CLK(clknet_leaf_68_clk),
    .D(net688),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14761_ (.CLK(clknet_leaf_68_clk),
    .D(net658),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14762_ (.CLK(clknet_leaf_24_clk),
    .D(net149),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14763_ (.CLK(clknet_leaf_24_clk),
    .D(net1458),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14764_ (.CLK(clknet_leaf_26_clk),
    .D(net1079),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14765_ (.CLK(clknet_leaf_21_clk),
    .D(net1450),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14766_ (.CLK(clknet_leaf_22_clk),
    .D(net381),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14767_ (.CLK(clknet_leaf_26_clk),
    .D(net1877),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14768_ (.CLK(clknet_leaf_69_clk),
    .D(net55),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _14769_ (.CLK(clknet_leaf_24_clk),
    .D(net1711),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _14770_ (.CLK(clknet_leaf_68_clk),
    .D(net445),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_1 _14771_ (.CLK(clknet_leaf_27_clk),
    .D(_00155_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _14772_ (.CLK(clknet_leaf_27_clk),
    .D(_00156_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14773_ (.CLK(clknet_leaf_33_clk),
    .D(_00157_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14774_ (.CLK(clknet_leaf_33_clk),
    .D(_00158_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14775_ (.CLK(clknet_leaf_27_clk),
    .D(net3447),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14776_ (.CLK(clknet_leaf_27_clk),
    .D(_00160_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14777_ (.CLK(clknet_leaf_27_clk),
    .D(_00161_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14778_ (.CLK(clknet_leaf_63_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14779_ (.CLK(clknet_leaf_67_clk),
    .D(net629),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14780_ (.CLK(clknet_leaf_67_clk),
    .D(net1418),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14781_ (.CLK(clknet_leaf_67_clk),
    .D(net2563),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14782_ (.CLK(clknet_leaf_14_clk),
    .D(_00002_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _14783_ (.CLK(clknet_leaf_34_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14784_ (.CLK(clknet_leaf_33_clk),
    .D(net2959),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14785_ (.CLK(clknet_leaf_34_clk),
    .D(net3020),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14786_ (.CLK(clknet_leaf_34_clk),
    .D(net3057),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14787_ (.CLK(clknet_leaf_33_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14788_ (.CLK(clknet_leaf_33_clk),
    .D(net3124),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14789_ (.CLK(clknet_leaf_34_clk),
    .D(net3047),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14790_ (.CLK(clknet_leaf_34_clk),
    .D(net3090),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14791_ (.CLK(clknet_leaf_33_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14792_ (.CLK(clknet_leaf_14_clk),
    .D(net887),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14793_ (.CLK(clknet_leaf_34_clk),
    .D(net946),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14794_ (.CLK(clknet_leaf_35_clk),
    .D(net2975),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14795_ (.CLK(clknet_leaf_26_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14796_ (.CLK(clknet_leaf_14_clk),
    .D(net559),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14797_ (.CLK(clknet_leaf_34_clk),
    .D(net2904),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14798_ (.CLK(clknet_leaf_34_clk),
    .D(net3073),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14799_ (.CLK(clknet_leaf_39_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[0] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14800_ (.CLK(clknet_leaf_39_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[1] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14801_ (.CLK(clknet_leaf_40_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[2] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14802_ (.CLK(clknet_leaf_39_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[3] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14803_ (.CLK(clknet_leaf_41_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[4] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14804_ (.CLK(clknet_leaf_41_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[5] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14805_ (.CLK(clknet_leaf_38_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[6] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14806_ (.CLK(clknet_leaf_38_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[7] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14807_ (.CLK(clknet_leaf_31_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[8] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14808_ (.CLK(clknet_leaf_31_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[9] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14809_ (.CLK(clknet_leaf_31_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[10] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14810_ (.CLK(clknet_leaf_31_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[11] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14811_ (.CLK(clknet_leaf_40_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[12] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14812_ (.CLK(clknet_leaf_39_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[13] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14813_ (.CLK(clknet_leaf_39_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[14] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14814_ (.CLK(clknet_leaf_39_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[15] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14815_ (.CLK(clknet_leaf_34_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[16] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14816_ (.CLK(clknet_leaf_32_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[17] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14817_ (.CLK(clknet_leaf_32_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[18] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14818_ (.CLK(clknet_leaf_41_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[19] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14819_ (.CLK(clknet_leaf_37_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[20] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14820_ (.CLK(clknet_leaf_37_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[21] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14821_ (.CLK(clknet_leaf_38_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[22] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14822_ (.CLK(clknet_leaf_38_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[23] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14823_ (.CLK(clknet_leaf_34_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[24] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14824_ (.CLK(clknet_leaf_31_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[25] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14825_ (.CLK(clknet_leaf_32_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[26] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14826_ (.CLK(clknet_leaf_41_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[27] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14827_ (.CLK(clknet_leaf_38_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[28] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14828_ (.CLK(clknet_leaf_37_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[29] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14829_ (.CLK(clknet_leaf_37_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[30] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14830_ (.CLK(clknet_leaf_37_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[31] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14831_ (.CLK(clknet_leaf_27_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[32] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14832_ (.CLK(clknet_leaf_28_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[33] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14833_ (.CLK(clknet_leaf_28_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[34] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14834_ (.CLK(clknet_leaf_25_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[35] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14835_ (.CLK(clknet_leaf_25_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[36] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14836_ (.CLK(clknet_leaf_25_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[37] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14837_ (.CLK(clknet_leaf_28_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[38] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14838_ (.CLK(clknet_leaf_28_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[39] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14839_ (.CLK(clknet_leaf_29_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[40] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14840_ (.CLK(clknet_leaf_27_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[41] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14841_ (.CLK(clknet_leaf_27_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[42] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14842_ (.CLK(clknet_leaf_29_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[43] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14843_ (.CLK(clknet_leaf_68_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[44] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14844_ (.CLK(clknet_leaf_68_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[45] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14845_ (.CLK(clknet_leaf_68_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.sr.ram_in[46] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14846_ (.CLK(clknet_leaf_40_clk),
    .D(net780),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14847_ (.CLK(clknet_leaf_39_clk),
    .D(net2227),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14848_ (.CLK(clknet_leaf_41_clk),
    .D(net274),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14849_ (.CLK(clknet_leaf_39_clk),
    .D(net2220),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14850_ (.CLK(clknet_leaf_41_clk),
    .D(net2749),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14851_ (.CLK(clknet_leaf_41_clk),
    .D(net1671),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14852_ (.CLK(clknet_leaf_41_clk),
    .D(net668),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14853_ (.CLK(clknet_leaf_38_clk),
    .D(net2226),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14854_ (.CLK(clknet_leaf_30_clk),
    .D(net256),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14855_ (.CLK(clknet_leaf_32_clk),
    .D(net2134),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14856_ (.CLK(clknet_leaf_31_clk),
    .D(net2802),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14857_ (.CLK(clknet_leaf_31_clk),
    .D(net1739),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14858_ (.CLK(clknet_leaf_39_clk),
    .D(net258),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14859_ (.CLK(clknet_leaf_39_clk),
    .D(net1858),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14860_ (.CLK(clknet_leaf_39_clk),
    .D(net2248),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14861_ (.CLK(clknet_leaf_39_clk),
    .D(net2107),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14862_ (.CLK(clknet_leaf_32_clk),
    .D(net683),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14863_ (.CLK(clknet_leaf_33_clk),
    .D(net205),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14864_ (.CLK(clknet_leaf_32_clk),
    .D(net972),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14865_ (.CLK(clknet_leaf_41_clk),
    .D(net1943),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14866_ (.CLK(clknet_leaf_37_clk),
    .D(net2037),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14867_ (.CLK(clknet_leaf_37_clk),
    .D(net2238),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14868_ (.CLK(clknet_leaf_38_clk),
    .D(net2027),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14869_ (.CLK(clknet_leaf_38_clk),
    .D(net2053),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14870_ (.CLK(clknet_leaf_34_clk),
    .D(net1724),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14871_ (.CLK(clknet_leaf_31_clk),
    .D(net2733),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14872_ (.CLK(clknet_leaf_32_clk),
    .D(net1319),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14873_ (.CLK(clknet_leaf_41_clk),
    .D(net2603),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14874_ (.CLK(clknet_leaf_37_clk),
    .D(net751),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14875_ (.CLK(clknet_leaf_37_clk),
    .D(net1534),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14876_ (.CLK(clknet_leaf_37_clk),
    .D(net2663),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14877_ (.CLK(clknet_leaf_37_clk),
    .D(net2041),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14878_ (.CLK(clknet_leaf_28_clk),
    .D(net220),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14879_ (.CLK(clknet_leaf_28_clk),
    .D(net2008),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14880_ (.CLK(clknet_leaf_28_clk),
    .D(net1900),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14881_ (.CLK(clknet_leaf_25_clk),
    .D(net2512),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14882_ (.CLK(clknet_leaf_25_clk),
    .D(net1631),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14883_ (.CLK(clknet_leaf_67_clk),
    .D(net561),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14884_ (.CLK(clknet_leaf_28_clk),
    .D(net1344),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14885_ (.CLK(clknet_leaf_28_clk),
    .D(net1308),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14886_ (.CLK(clknet_leaf_29_clk),
    .D(net1784),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14887_ (.CLK(clknet_leaf_27_clk),
    .D(net1171),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14888_ (.CLK(clknet_leaf_27_clk),
    .D(net842),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14889_ (.CLK(clknet_leaf_29_clk),
    .D(net2217),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14890_ (.CLK(clknet_leaf_68_clk),
    .D(net2798),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14891_ (.CLK(clknet_leaf_68_clk),
    .D(net1202),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14892_ (.CLK(clknet_leaf_68_clk),
    .D(net2665),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14893_ (.CLK(clknet_leaf_40_clk),
    .D(net1479),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14894_ (.CLK(clknet_leaf_39_clk),
    .D(net1707),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14895_ (.CLK(clknet_leaf_41_clk),
    .D(net2490),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14896_ (.CLK(clknet_leaf_39_clk),
    .D(net1488),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14897_ (.CLK(clknet_leaf_41_clk),
    .D(net1323),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14898_ (.CLK(clknet_leaf_41_clk),
    .D(net2764),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14899_ (.CLK(clknet_leaf_41_clk),
    .D(net2421),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14900_ (.CLK(clknet_leaf_38_clk),
    .D(net2451),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14901_ (.CLK(clknet_leaf_31_clk),
    .D(net108),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14902_ (.CLK(clknet_leaf_31_clk),
    .D(net206),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14903_ (.CLK(clknet_leaf_31_clk),
    .D(net1856),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14904_ (.CLK(clknet_leaf_31_clk),
    .D(net1740),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14905_ (.CLK(clknet_leaf_40_clk),
    .D(net777),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14906_ (.CLK(clknet_leaf_39_clk),
    .D(net1456),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14907_ (.CLK(clknet_leaf_39_clk),
    .D(net2767),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14908_ (.CLK(clknet_leaf_39_clk),
    .D(net1270),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14909_ (.CLK(clknet_leaf_32_clk),
    .D(net881),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14910_ (.CLK(clknet_leaf_32_clk),
    .D(net1709),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14911_ (.CLK(clknet_leaf_32_clk),
    .D(net870),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14912_ (.CLK(clknet_leaf_42_clk),
    .D(net759),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14913_ (.CLK(clknet_leaf_37_clk),
    .D(net1513),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14914_ (.CLK(clknet_leaf_37_clk),
    .D(net1522),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14915_ (.CLK(clknet_leaf_38_clk),
    .D(net2592),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14916_ (.CLK(clknet_leaf_38_clk),
    .D(net1793),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14917_ (.CLK(clknet_leaf_34_clk),
    .D(net1031),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14918_ (.CLK(clknet_leaf_31_clk),
    .D(net2469),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14919_ (.CLK(clknet_leaf_31_clk),
    .D(net204),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14920_ (.CLK(clknet_leaf_42_clk),
    .D(net745),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14921_ (.CLK(clknet_leaf_38_clk),
    .D(net396),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14922_ (.CLK(clknet_leaf_37_clk),
    .D(net1633),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14923_ (.CLK(clknet_leaf_37_clk),
    .D(net1204),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14924_ (.CLK(clknet_leaf_37_clk),
    .D(net1196),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14925_ (.CLK(clknet_leaf_28_clk),
    .D(net2022),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _14926_ (.CLK(clknet_leaf_28_clk),
    .D(net2778),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _14927_ (.CLK(clknet_leaf_28_clk),
    .D(net1667),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _14928_ (.CLK(clknet_leaf_25_clk),
    .D(net2857),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _14929_ (.CLK(clknet_leaf_25_clk),
    .D(net2275),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _14930_ (.CLK(clknet_leaf_67_clk),
    .D(net2633),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _14931_ (.CLK(clknet_leaf_28_clk),
    .D(net1803),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _14932_ (.CLK(clknet_leaf_25_clk),
    .D(net448),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _14933_ (.CLK(clknet_leaf_29_clk),
    .D(net2343),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _14934_ (.CLK(clknet_leaf_28_clk),
    .D(net210),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _14935_ (.CLK(clknet_leaf_27_clk),
    .D(net850),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _14936_ (.CLK(clknet_leaf_29_clk),
    .D(net2310),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _14937_ (.CLK(clknet_leaf_68_clk),
    .D(net1806),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _14938_ (.CLK(clknet_leaf_68_clk),
    .D(net1596),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _14939_ (.CLK(clknet_leaf_68_clk),
    .D(net1928),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _14940_ (.CLK(clknet_leaf_40_clk),
    .D(net922),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14941_ (.CLK(clknet_leaf_39_clk),
    .D(net1291),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14942_ (.CLK(clknet_leaf_41_clk),
    .D(net2862),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14943_ (.CLK(clknet_leaf_39_clk),
    .D(net1302),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14944_ (.CLK(clknet_leaf_41_clk),
    .D(net2476),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14945_ (.CLK(clknet_leaf_42_clk),
    .D(net735),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14946_ (.CLK(clknet_leaf_41_clk),
    .D(net2229),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14947_ (.CLK(clknet_leaf_41_clk),
    .D(net654),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14948_ (.CLK(clknet_leaf_31_clk),
    .D(net2406),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14949_ (.CLK(clknet_leaf_31_clk),
    .D(net1446),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14950_ (.CLK(clknet_leaf_29_clk),
    .D(net249),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14951_ (.CLK(clknet_leaf_29_clk),
    .D(net243),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14952_ (.CLK(clknet_leaf_38_clk),
    .D(net257),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14953_ (.CLK(clknet_leaf_39_clk),
    .D(net2652),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14954_ (.CLK(clknet_leaf_39_clk),
    .D(net1224),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14955_ (.CLK(clknet_leaf_38_clk),
    .D(net418),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14956_ (.CLK(clknet_leaf_32_clk),
    .D(net879),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14957_ (.CLK(clknet_leaf_33_clk),
    .D(net207),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14958_ (.CLK(clknet_leaf_32_clk),
    .D(net886),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14959_ (.CLK(clknet_leaf_31_clk),
    .D(net288),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14960_ (.CLK(clknet_leaf_38_clk),
    .D(net300),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14961_ (.CLK(clknet_leaf_38_clk),
    .D(net420),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14962_ (.CLK(clknet_leaf_38_clk),
    .D(net1543),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14963_ (.CLK(clknet_leaf_38_clk),
    .D(net1482),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14964_ (.CLK(clknet_leaf_32_clk),
    .D(net662),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14965_ (.CLK(clknet_leaf_31_clk),
    .D(net1738),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14966_ (.CLK(clknet_leaf_31_clk),
    .D(net2178),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14967_ (.CLK(clknet_leaf_41_clk),
    .D(net320),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14968_ (.CLK(clknet_leaf_38_clk),
    .D(net1315),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14969_ (.CLK(clknet_leaf_37_clk),
    .D(net1214),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14970_ (.CLK(clknet_leaf_37_clk),
    .D(net1742),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14971_ (.CLK(clknet_leaf_38_clk),
    .D(net405),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14972_ (.CLK(clknet_leaf_25_clk),
    .D(net393),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14973_ (.CLK(clknet_leaf_25_clk),
    .D(net422),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14974_ (.CLK(clknet_leaf_28_clk),
    .D(net1939),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14975_ (.CLK(clknet_leaf_25_clk),
    .D(net1552),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14976_ (.CLK(clknet_leaf_67_clk),
    .D(net626),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14977_ (.CLK(clknet_leaf_67_clk),
    .D(net2198),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14978_ (.CLK(clknet_leaf_28_clk),
    .D(net2697),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14979_ (.CLK(clknet_leaf_67_clk),
    .D(net608),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14980_ (.CLK(clknet_leaf_28_clk),
    .D(net500),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14981_ (.CLK(clknet_leaf_28_clk),
    .D(net1306),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14982_ (.CLK(clknet_leaf_27_clk),
    .D(net930),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14983_ (.CLK(clknet_leaf_29_clk),
    .D(net2588),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14984_ (.CLK(clknet_leaf_69_clk),
    .D(net63),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fd ));
 sky130_fd_sc_hd__dfxtp_1 _14985_ (.CLK(clknet_leaf_69_clk),
    .D(net59),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fds ));
 sky130_fd_sc_hd__dfxtp_1 _14986_ (.CLK(clknet_leaf_69_clk),
    .D(net61),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fde ));
 sky130_fd_sc_hd__dfxtp_2 _14987_ (.CLK(clknet_leaf_27_clk),
    .D(_00162_),
    .Q(\c.genblk1.genblk1.subs.c0.cfgd ));
 sky130_fd_sc_hd__dfxtp_1 _14988_ (.CLK(clknet_leaf_27_clk),
    .D(_00163_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14989_ (.CLK(clknet_leaf_27_clk),
    .D(_00164_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14990_ (.CLK(clknet_leaf_33_clk),
    .D(net3276),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14991_ (.CLK(clknet_leaf_33_clk),
    .D(_00166_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14992_ (.CLK(clknet_leaf_33_clk),
    .D(_00167_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14993_ (.CLK(clknet_leaf_33_clk),
    .D(_00168_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14994_ (.CLK(clknet_leaf_24_clk),
    .D(_00169_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ));
 sky130_fd_sc_hd__dfxtp_1 _14995_ (.CLK(clknet_leaf_63_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14996_ (.CLK(clknet_leaf_67_clk),
    .D(net541),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14997_ (.CLK(clknet_leaf_68_clk),
    .D(net526),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14998_ (.CLK(clknet_leaf_68_clk),
    .D(net1463),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14999_ (.CLK(clknet_leaf_34_clk),
    .D(_00003_),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.half_q ));
 sky130_fd_sc_hd__dfxtp_1 _15000_ (.CLK(clknet_leaf_34_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15001_ (.CLK(clknet_leaf_35_clk),
    .D(net2958),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15002_ (.CLK(clknet_leaf_38_clk),
    .D(net2964),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15003_ (.CLK(clknet_leaf_38_clk),
    .D(net3083),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15004_ (.CLK(clknet_leaf_34_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[1] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15005_ (.CLK(clknet_leaf_35_clk),
    .D(net2961),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15006_ (.CLK(clknet_leaf_35_clk),
    .D(net3045),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15007_ (.CLK(clknet_leaf_35_clk),
    .D(net3079),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15008_ (.CLK(clknet_leaf_41_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[2] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15009_ (.CLK(clknet_leaf_38_clk),
    .D(net2967),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15010_ (.CLK(clknet_leaf_41_clk),
    .D(net2987),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15011_ (.CLK(clknet_leaf_38_clk),
    .D(net2972),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15012_ (.CLK(clknet_leaf_32_clk),
    .D(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[3] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15013_ (.CLK(clknet_leaf_32_clk),
    .D(net3116),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15014_ (.CLK(clknet_leaf_32_clk),
    .D(net3123),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15015_ (.CLK(clknet_leaf_38_clk),
    .D(net2965),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15016_ (.CLK(clknet_leaf_65_clk),
    .D(net3417),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__dfxtp_4 _15017_ (.CLK(clknet_leaf_65_clk),
    .D(net3490),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15018_ (.CLK(clknet_leaf_66_clk),
    .D(net3665),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15019_ (.CLK(clknet_leaf_66_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[3] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15020_ (.CLK(clknet_leaf_72_clk),
    .D(net3392),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15021_ (.CLK(clknet_leaf_66_clk),
    .D(net3495),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15022_ (.CLK(clknet_leaf_63_clk),
    .D(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[6] ),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15023_ (.CLK(clknet_leaf_65_clk),
    .D(net3633),
    .Q(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(cfg),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(net51),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(net43),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(net42),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(net54),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(net44),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(net37),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(net39),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(net50),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(net76),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(up_i[0]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(up_i[10]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(up_i[11]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(up_i[12]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(up_i[13]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(up_i[14]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(up_i[15]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(up_i[1]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(up_i[2]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(up_i[3]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(up_i[4]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(up_i[5]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(up_i[6]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(up_i[7]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(up_i[8]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(up_i[9]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(cfgd));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(up_o[0]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(up_o[1]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(up_o[2]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(up_o[3]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(up_o[4]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(up_o[5]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(up_o[6]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(up_o[7]));
 sky130_fd_sc_hd__conb_1 x64_36 (.LO(net36));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_opt_2_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_opt_3_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_opt_1_0_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_clk (.A(clknet_1_0_0_clk),
    .X(clknet_1_0_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_clk (.A(clknet_1_1_0_clk),
    .X(clknet_1_1_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_opt_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_opt_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_opt_3_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(grst),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net7),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(m[0]),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net8),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net4215),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(cfg_i[2]),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(cfg_i[1]),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(cfg_i[4]),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][20] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][31] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][19] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][23] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][16] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(m[1]),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(cfg_i[0]),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][23] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][39] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(cfg_i[3]),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][27] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][7] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][31] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(rst),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][17] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][32] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][0] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][36] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][11] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][25] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][27] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][10] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][34] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][30] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][36] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][38] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][38] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][23] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][37] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][35] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\c.genblk1.genblk1.subs.sw.up.x.o[4] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\c.cfg_i_q[4] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\c.genblk1.genblk1.subs.sw.up.x.o[7] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][0] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[23] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\c.genblk1.genblk1.subs.sw.up.x.o_[5] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][1] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][37] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][20] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][34] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][18] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][39] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][35] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][2] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][14] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][22] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][35] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][17] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][23] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][9] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][38] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][0] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][30] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][27] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][33] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][26] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][2] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][23] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][11] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][29] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][12] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][14] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][10] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][28] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][0] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][26] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][23] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][21] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][19] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][6] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][17] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][23] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][17] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][16] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][20] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][24] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][18] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][25] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][25] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][3] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][20] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][9] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][11] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][15] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][34] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][26] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][31] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][6] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][26] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][32] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][15] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][27] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][32] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][1] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][7] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][32] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][31] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][15] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][2] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][33] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][0] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][16] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][14] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][13] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][16] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][21] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][38] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][17] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][10] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][2] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][27] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][37] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][9] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][39] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][18] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][1] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][24] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][26] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][10] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][11] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][6] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][5] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][39] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][21] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][1] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][2] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][30] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][12] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][9] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][13] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][29] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][5] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][14] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][36] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][12] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][7] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][29] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][16] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][27] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][36] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][3] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][1] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][29] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][3] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][31] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][2] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][10] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][39] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][33] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][31] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][30] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][2] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][5] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\c.genblk1.genblk1.subs.c0.m[0] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][28] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][17] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][31] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][0] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][24] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][10] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][23] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][35] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][37] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][1] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][39] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][22] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][8] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][36] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][8] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][31] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][15] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][38] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][22] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][15] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][37] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][8] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][8] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][20] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][4] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][39] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\c.genblk1.genblk1.subs.c0.grst ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][23] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][18] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][1] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][31] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\c.genblk1.genblk1.subs.sw.up.x.o[3] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][20] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][6] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][18] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][20] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][4] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][17] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][16] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][38] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][21] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][39] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][30] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][37] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][19] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][22] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][12] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][7] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][14] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][39] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][26] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][7] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][21] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][30] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][16] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][36] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][19] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][23] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][0] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][31] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][30] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][1] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][17] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][10] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][39] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\c.cfg_i_q[3] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][16] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][18] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][22] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][11] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][30] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][10] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][36] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][29] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][33] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][36] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][22] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][21] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][16] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][20] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][20] ),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][22] ),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][0] ),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][35] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][15] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][15] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][35] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][24] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][35] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][38] ),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][5] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][0] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][6] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][16] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][22] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][18] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][17] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][30] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][4] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][17] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][20] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][10] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][10] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][31] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][22] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][8] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][21] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][3] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][13] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][34] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][21] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][14] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][1] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][32] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][28] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][29] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][33] ),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][18] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][11] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][5] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][28] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][30] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[0] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][5] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][13] ),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][6] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][4] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][24] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][4] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][18] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][9] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][20] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][5] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][8] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][3] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][17] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][40] ),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][16] ),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][12] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][23] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\c.genblk1.genblk1.subs.c0.rst ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][4] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][16] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][30] ),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][19] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][23] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][7] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][37] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][9] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][20] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][22] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][26] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][19] ),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][24] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][26] ),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][29] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][7] ),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][23] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][4] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][13] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][0] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][18] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][8] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][11] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][28] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][11] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][13] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][27] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][33] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][10] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][7] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][37] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][1] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][24] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][27] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][14] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][42] ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][3] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][9] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][16] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][7] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][25] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][27] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][18] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][15] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][15] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][36] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][11] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][27] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][4] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][12] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][1] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][11] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][41] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][1] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(\c.cfg_i_q[1] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][4] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][19] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][25] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][24] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][20] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][36] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][38] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][22] ),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][9] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][14] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][36] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][1] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][24] ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][25] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][34] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][19] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][37] ),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][2] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][31] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(\c.cfg_i_q[0] ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][6] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][11] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][24] ),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][4] ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][7] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][1] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][11] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][28] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][34] ),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][14] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][35] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][39] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][1] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][17] ),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][19] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][32] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][44] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][16] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][15] ),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][38] ),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][18] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][4] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][0] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][0] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][32] ),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][3] ),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][2] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][14] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(\c.genblk1.genblk1.subs.c0.m[1] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][25] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][16] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][15] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][10] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][1] ),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][7] ),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][16] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][25] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][14] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][2] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][34] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][37] ),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][11] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][5] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][16] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][1] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][39] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][30] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][27] ),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][38] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][29] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][6] ),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][38] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][8] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][12] ),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][38] ),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][24] ),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][19] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][11] ),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][31] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][37] ),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][7] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][0] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][13] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][34] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][28] ),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][8] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][29] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][5] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][13] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][27] ),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][4] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][33] ),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][6] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][36] ),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][28] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][16] ),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][18] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][45] ),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][36] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[1] ),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][25] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][11] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][30] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][38] ),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][14] ),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][21] ),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][45] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][39] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][32] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][5] ),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][16] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][29] ),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][8] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][6] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][2] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][39] ),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][5] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][18] ),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][18] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][11] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][40] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][37] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][40] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][2] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][15] ),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][35] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][29] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][18] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][1] ),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[0] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][10] ),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][17] ),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][16] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][35] ),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][12] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][21] ),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][21] ),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][3] ),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1794 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][15] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][26] ),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][24] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][39] ),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][29] ),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][8] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][12] ),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][23] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1808 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][27] ),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][7] ),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][26] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][16] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1827 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][33] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1831 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][14] ),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1835 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][19] ),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][29] ),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][2] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][21] ),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][35] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][11] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][44] ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1849 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1850 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1851 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][25] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1852 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1853 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1854 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1855 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][37] ),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1856 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][3] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1857 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1858 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1859 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][29] ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1860 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][4] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1861 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1862 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1863 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][26] ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1864 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1865 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][28] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1866 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1867 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][36] ),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1868 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1869 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1870 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1871 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][15] ),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1872 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][26] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1873 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1874 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1875 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][37] ),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1876 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][13] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1877 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][2] ),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1878 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1879 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1880 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][8] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1881 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][14] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1882 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1883 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1884 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][20] ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1885 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1886 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1887 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][32] ),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1888 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1889 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1890 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][24] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1891 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1892 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][46] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1893 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][17] ),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1894 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1895 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1896 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][20] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1897 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][29] ),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1898 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][23] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1899 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1900 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1901 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][7] ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1902 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][33] ),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1903 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1904 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1905 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1906 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1907 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1908 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][9] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1909 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1910 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1911 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1912 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][33] ),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1913 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][25] ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1914 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1915 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1916 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1917 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][37] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1918 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1919 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1920 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1921 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1922 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1923 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1924 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1925 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1926 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][42] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1927 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1928 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1929 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][18] ),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1930 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][19] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1931 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1932 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][31] ),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1933 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1934 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][21] ),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1935 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1936 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][27] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1937 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1938 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1939 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1940 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1941 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][19] ),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1942 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1943 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][31] ),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1944 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1945 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][31] ),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1946 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1947 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1948 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][21] ),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1949 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1950 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][12] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1951 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1952 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1953 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][13] ),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1954 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1955 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][2] ),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1956 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][35] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1957 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1958 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1959 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][10] ),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1960 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1961 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1962 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][15] ),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1963 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1964 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1965 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][9] ),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1966 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1967 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][29] ),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1968 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1969 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1970 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][25] ),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1971 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][26] ),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1972 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1973 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][34] ),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1974 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][6] ),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1975 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1976 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1977 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1978 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][3] ),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1979 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1980 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1981 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][30] ),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1982 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1983 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1984 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][18] ),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1985 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][33] ),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1986 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1987 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1988 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1989 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][2] ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1990 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1991 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][22] ),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1992 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][9] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1993 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][25] ),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1994 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1995 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1996 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1997 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][41] ),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1998 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][2] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1999 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2000 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2001 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2002 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2003 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2004 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][21] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2005 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2006 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2007 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2008 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][34] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2009 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][19] ),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2010 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][3] ),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2011 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2012 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2013 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][11] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2014 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][35] ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2015 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2016 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][4] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2017 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2018 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2019 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2020 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2021 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][10] ),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2022 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2023 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2024 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2025 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2026 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][21] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2027 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][25] ),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2028 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2029 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2030 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2031 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][19] ),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2032 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][33] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2033 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][18] ),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2034 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2035 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2036 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2037 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][34] ),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2038 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][32] ),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2039 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2040 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][39] ),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2041 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2042 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.qs[2] ),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2043 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2044 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2045 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2046 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][31] ),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2047 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2048 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2049 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2050 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2051 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][31] ),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2052 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2053 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2054 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2055 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2056 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2057 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][43] ),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2058 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][3] ),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2059 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2060 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][34] ),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2061 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][39] ),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2062 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][35] ),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2063 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][42] ),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2064 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2065 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2066 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2067 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2068 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][20] ),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2069 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2070 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][20] ),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2071 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2072 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2073 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][33] ),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2074 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][36] ),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2075 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2076 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2077 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2078 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][33] ),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2079 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2080 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][26] ),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2081 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][40] ),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2082 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][6] ),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2083 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2084 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2085 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2086 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][27] ),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2087 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2088 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][19] ),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2089 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2090 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][23] ),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2091 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2092 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][37] ),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2093 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][22] ),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2094 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][28] ),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2095 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][22] ),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2096 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][30] ),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2097 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][32] ),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2098 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2099 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2100 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2101 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2102 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][9] ),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2103 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2104 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][38] ),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2105 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2106 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][24] ),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2107 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][13] ),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2108 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][22] ),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2109 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2110 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2111 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][9] ),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2112 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][1] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2113 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2114 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][7] ),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2115 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2116 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][19] ),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2117 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2118 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][10] ),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2119 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][12] ),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2120 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2121 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2122 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2123 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2124 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][33] ),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2125 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][17] ),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2126 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2127 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][8] ),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2128 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2129 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][29] ),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2130 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][25] ),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2131 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][6] ),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2132 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][23] ),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2133 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2134 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2135 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2136 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2137 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][6] ),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2138 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][32] ),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2139 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][15] ),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2140 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2141 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2142 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][26] ),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2143 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2144 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2145 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2146 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2147 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][4] ),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2148 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2149 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2150 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2151 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][34] ),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2152 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][19] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2153 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2154 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2155 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2156 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][15] ),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2157 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2158 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][15] ),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2159 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][3] ),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2160 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][8] ),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2161 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ),
    .X(net2197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2162 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][37] ),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2163 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2164 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2165 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2166 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2167 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2168 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][5] ),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2169 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][25] ),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2170 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2171 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][28] ),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2172 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2173 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][2] ),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2174 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][46] ),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2175 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2176 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][12] ),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2177 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][27] ),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2178 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2179 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[2] ),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2180 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2181 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][43] ),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2182 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][4] ),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2183 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][26] ),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2184 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2185 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2186 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2187 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2188 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][36] ),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2189 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2190 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2191 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2192 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][12] ),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2193 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][6] ),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2194 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][46] ),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2195 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][24] ),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2196 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2197 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2198 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2199 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2200 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2201 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2202 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2203 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][45] ),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2204 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2205 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][7] ),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2206 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][19] ),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2207 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2208 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2209 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2210 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][25] ),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2211 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][20] ),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2212 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2213 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2214 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2215 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][12] ),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2216 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2217 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][21] ),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2218 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2219 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][35] ),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2220 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2221 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][10] ),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2222 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][6] ),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2223 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2224 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][27] ),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2225 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2226 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2227 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2228 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][18] ),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2229 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2230 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][21] ),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2231 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][4] ),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2232 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][43] ),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2233 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2234 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2235 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2236 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2237 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2238 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2239 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2240 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][8] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2241 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2242 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2243 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2244 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2245 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][10] ),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2246 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2247 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2248 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2249 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2250 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][34] ),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2251 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][3] ),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2252 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2253 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2254 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2255 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2256 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2257 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2258 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2259 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2260 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][23] ),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2261 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2262 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][5] ),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2263 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2264 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2265 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2266 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2267 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][27] ),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2268 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2269 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][37] ),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2270 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2271 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2272 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2273 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][27] ),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2274 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2275 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2276 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][15] ),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2277 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2278 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2279 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2280 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2281 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][42] ),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2282 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2283 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2284 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][19] ),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2285 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][42] ),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2286 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2287 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2288 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][32] ),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2289 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[1] ),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2290 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][28] ),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2291 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2292 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][14] ),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2293 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][0] ),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2294 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2295 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2296 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][24] ),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2297 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][46] ),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2298 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2299 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][22] ),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2300 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][32] ),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2301 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][24] ),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2302 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2303 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][34] ),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2304 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2305 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][43] ),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2306 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][10] ),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2307 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2308 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][39] ),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2309 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][8] ),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2310 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][28] ),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2311 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2312 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2313 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][8] ),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2314 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2315 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2316 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2317 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][36] ),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2318 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2319 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][9] ),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2320 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][26] ),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2321 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][4] ),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2322 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][3] ),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2323 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2324 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2325 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2326 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][8] ),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2327 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2328 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][29] ),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2329 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2330 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2331 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][25] ),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2332 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2333 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][1] ),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2334 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2335 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2336 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][3] ),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2337 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2338 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][5] ),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2339 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][8] ),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2340 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][44] ),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2341 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][5] ),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2342 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][0] ),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2343 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][7] ),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2344 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][45] ),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2345 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2346 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][15] ),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2347 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2348 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2349 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][6] ),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2350 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[2] ),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2351 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2352 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][18] ),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2353 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2354 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][45] ),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2355 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2356 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][14] ),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2357 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ),
    .X(net2393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2358 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][45] ),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2359 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2360 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2361 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][6] ),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2362 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][33] ),
    .X(net2398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2363 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[1] ),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2364 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ),
    .X(net2400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2365 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][6] ),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2366 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2367 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2368 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2369 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][7] ),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2370 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][8] ),
    .X(net2406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2371 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][45] ),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2372 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][1] ),
    .X(net2408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2373 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][14] ),
    .X(net2409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2374 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][3] ),
    .X(net2410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2375 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ),
    .X(net2411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2376 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][43] ),
    .X(net2412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2377 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][22] ),
    .X(net2413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2378 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ),
    .X(net2414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2379 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][22] ),
    .X(net2415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2380 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ),
    .X(net2416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2381 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][39] ),
    .X(net2417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2382 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][25] ),
    .X(net2418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2383 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][36] ),
    .X(net2419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2384 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][44] ),
    .X(net2420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2385 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][6] ),
    .X(net2421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2386 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][21] ),
    .X(net2422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2387 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][26] ),
    .X(net2423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2388 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][29] ),
    .X(net2424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2389 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][17] ),
    .X(net2425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2390 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][8] ),
    .X(net2426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2391 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][20] ),
    .X(net2427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2392 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ),
    .X(net2428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2393 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ),
    .X(net2429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2394 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ),
    .X(net2430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2395 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][24] ),
    .X(net2431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2396 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][7] ),
    .X(net2432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2397 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ),
    .X(net2433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2398 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ),
    .X(net2434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2399 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][23] ),
    .X(net2435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2400 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][9] ),
    .X(net2436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2401 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ),
    .X(net2437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2402 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][21] ),
    .X(net2438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2403 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][13] ),
    .X(net2439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2404 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][12] ),
    .X(net2440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2405 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ),
    .X(net2441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2406 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][45] ),
    .X(net2442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2407 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ),
    .X(net2443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2408 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ),
    .X(net2444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2409 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][33] ),
    .X(net2445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2410 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ),
    .X(net2446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2411 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][40] ),
    .X(net2447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2412 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][3] ),
    .X(net2448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2413 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][43] ),
    .X(net2449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2414 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ),
    .X(net2450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2415 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ),
    .X(net2451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2416 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][0] ),
    .X(net2452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2417 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][11] ),
    .X(net2453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2418 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ),
    .X(net2454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2419 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][43] ),
    .X(net2455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2420 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ),
    .X(net2456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2421 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ),
    .X(net2457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2422 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][45] ),
    .X(net2458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2423 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ),
    .X(net2459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2424 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ),
    .X(net2460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2425 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ),
    .X(net2461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2426 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ),
    .X(net2462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2427 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][25] ),
    .X(net2463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2428 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][11] ),
    .X(net2464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2429 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ),
    .X(net2465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2430 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][35] ),
    .X(net2466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2431 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][9] ),
    .X(net2467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2432 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][16] ),
    .X(net2468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2433 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][25] ),
    .X(net2469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2434 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][11] ),
    .X(net2470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2435 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ),
    .X(net2471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2436 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][22] ),
    .X(net2472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2437 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][10] ),
    .X(net2473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2438 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][17] ),
    .X(net2474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2439 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][45] ),
    .X(net2475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2440 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ),
    .X(net2476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2441 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ),
    .X(net2477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2442 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ),
    .X(net2478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2443 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][16] ),
    .X(net2479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2444 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][34] ),
    .X(net2480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2445 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][30] ),
    .X(net2481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2446 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ),
    .X(net2482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2447 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ),
    .X(net2483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2448 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][13] ),
    .X(net2484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2449 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][32] ),
    .X(net2485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2450 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][40] ),
    .X(net2486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2451 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][0] ),
    .X(net2487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2452 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][15] ),
    .X(net2488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2453 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ),
    .X(net2489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2454 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ),
    .X(net2490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2455 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][11] ),
    .X(net2491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2456 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ),
    .X(net2492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2457 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][28] ),
    .X(net2493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2458 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][41] ),
    .X(net2494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2459 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][36] ),
    .X(net2495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2460 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][0] ),
    .X(net2496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2461 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][0] ),
    .X(net2497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2462 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ),
    .X(net2498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2463 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ),
    .X(net2499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2464 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][12] ),
    .X(net2500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2465 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][3] ),
    .X(net2501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2466 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][13] ),
    .X(net2502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2467 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ),
    .X(net2503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2468 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ),
    .X(net2504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2469 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][5] ),
    .X(net2505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2470 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ),
    .X(net2506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2471 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][13] ),
    .X(net2507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2472 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][5] ),
    .X(net2508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2473 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][37] ),
    .X(net2509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2474 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][41] ),
    .X(net2510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2475 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][12] ),
    .X(net2511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2476 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][35] ),
    .X(net2512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2477 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ),
    .X(net2513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2478 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][31] ),
    .X(net2514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2479 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ),
    .X(net2515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2480 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ),
    .X(net2516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2481 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ),
    .X(net2517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2482 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ),
    .X(net2518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2483 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][32] ),
    .X(net2519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2484 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ),
    .X(net2520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2485 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ),
    .X(net2521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2486 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ),
    .X(net2522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2487 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][11] ),
    .X(net2523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2488 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][28] ),
    .X(net2524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2489 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][23] ),
    .X(net2525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2490 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ),
    .X(net2526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2491 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][44] ),
    .X(net2527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2492 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][36] ),
    .X(net2528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2493 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][17] ),
    .X(net2529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2494 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][28] ),
    .X(net2530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2495 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ),
    .X(net2531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2496 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][5] ),
    .X(net2532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2497 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][38] ),
    .X(net2533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2498 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ),
    .X(net2534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2499 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][23] ),
    .X(net2535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2500 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][32] ),
    .X(net2536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2501 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][27] ),
    .X(net2537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2502 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ),
    .X(net2538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2503 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ),
    .X(net2539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2504 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ),
    .X(net2540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2505 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ),
    .X(net2541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2506 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][19] ),
    .X(net2542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2507 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][14] ),
    .X(net2543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2508 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ),
    .X(net2544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2509 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ),
    .X(net2545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2510 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.qs[0] ),
    .X(net2546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2511 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][29] ),
    .X(net2547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2512 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][18] ),
    .X(net2548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2513 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ),
    .X(net2549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2514 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][9] ),
    .X(net2550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2515 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][31] ),
    .X(net2551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2516 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][8] ),
    .X(net2552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2517 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ),
    .X(net2553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2518 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][36] ),
    .X(net2554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2519 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][27] ),
    .X(net2555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2520 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][39] ),
    .X(net2556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2521 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][26] ),
    .X(net2557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2522 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ),
    .X(net2558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2523 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ),
    .X(net2559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2524 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ),
    .X(net2560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2525 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ),
    .X(net2561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2526 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][5] ),
    .X(net2562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2527 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.qs[2] ),
    .X(net2563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2528 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][17] ),
    .X(net2564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2529 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][27] ),
    .X(net2565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2530 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][17] ),
    .X(net2566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2531 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][35] ),
    .X(net2567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2532 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][43] ),
    .X(net2568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2533 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][44] ),
    .X(net2569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2534 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][24] ),
    .X(net2570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2535 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][7] ),
    .X(net2571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2536 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][2] ),
    .X(net2572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2537 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ),
    .X(net2573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2538 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][18] ),
    .X(net2574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2539 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][24] ),
    .X(net2575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2540 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ),
    .X(net2576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2541 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][24] ),
    .X(net2577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2542 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ),
    .X(net2578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2543 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][14] ),
    .X(net2579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2544 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ),
    .X(net2580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2545 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][13] ),
    .X(net2581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2546 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][31] ),
    .X(net2582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2547 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ),
    .X(net2583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2548 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ),
    .X(net2584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2549 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][20] ),
    .X(net2585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2550 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][5] ),
    .X(net2586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2551 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][4] ),
    .X(net2587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2552 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ),
    .X(net2588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2553 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][33] ),
    .X(net2589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2554 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][35] ),
    .X(net2590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2555 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ),
    .X(net2591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2556 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][22] ),
    .X(net2592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2557 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ),
    .X(net2593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2558 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][13] ),
    .X(net2594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2559 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][13] ),
    .X(net2595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2560 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][9] ),
    .X(net2596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2561 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][4] ),
    .X(net2597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2562 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ),
    .X(net2598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2563 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ),
    .X(net2599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2564 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][41] ),
    .X(net2600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2565 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][14] ),
    .X(net2601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2566 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][13] ),
    .X(net2602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2567 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][27] ),
    .X(net2603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2568 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][22] ),
    .X(net2604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2569 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][12] ),
    .X(net2605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2570 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][38] ),
    .X(net2606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2571 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ),
    .X(net2607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2572 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][2] ),
    .X(net2608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2573 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ),
    .X(net2609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2574 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[2][38] ),
    .X(net2610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2575 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][6] ),
    .X(net2611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2576 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][13] ),
    .X(net2612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2577 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][2] ),
    .X(net2613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2578 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][24] ),
    .X(net2614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2579 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][44] ),
    .X(net2615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2580 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ),
    .X(net2616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2581 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][42] ),
    .X(net2617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2582 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ),
    .X(net2618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2583 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][42] ),
    .X(net2619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2584 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.qs[0] ),
    .X(net2620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2585 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][8] ),
    .X(net2621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2586 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][4] ),
    .X(net2622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2587 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][9] ),
    .X(net2623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2588 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][19] ),
    .X(net2624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2589 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][2] ),
    .X(net2625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2590 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][31] ),
    .X(net2626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2591 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][12] ),
    .X(net2627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2592 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.qs[1] ),
    .X(net2628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2593 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][33] ),
    .X(net2629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2594 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][9] ),
    .X(net2630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2595 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][10] ),
    .X(net2631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2596 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][6] ),
    .X(net2632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2597 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][37] ),
    .X(net2633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2598 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][24] ),
    .X(net2634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2599 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ),
    .X(net2635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2600 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][45] ),
    .X(net2636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2601 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ),
    .X(net2637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2602 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][32] ),
    .X(net2638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2603 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][34] ),
    .X(net2639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2604 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][3] ),
    .X(net2640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2605 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][44] ),
    .X(net2641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2606 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][7] ),
    .X(net2642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2607 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ),
    .X(net2643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2608 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ),
    .X(net2644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2609 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ),
    .X(net2645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2610 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ),
    .X(net2646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2611 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][10] ),
    .X(net2647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2612 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][18] ),
    .X(net2648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2613 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][11] ),
    .X(net2649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2614 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][0] ),
    .X(net2650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2615 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ),
    .X(net2651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2616 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ),
    .X(net2652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2617 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][10] ),
    .X(net2653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2618 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][26] ),
    .X(net2654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2619 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][17] ),
    .X(net2655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2620 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ),
    .X(net2656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2621 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ),
    .X(net2657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2622 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][10] ),
    .X(net2658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2623 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][42] ),
    .X(net2659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2624 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][33] ),
    .X(net2660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2625 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][6] ),
    .X(net2661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2626 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][35] ),
    .X(net2662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2627 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][30] ),
    .X(net2663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2628 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][19] ),
    .X(net2664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2629 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][46] ),
    .X(net2665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2630 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][20] ),
    .X(net2666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2631 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][12] ),
    .X(net2667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2632 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][5] ),
    .X(net2668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2633 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][15] ),
    .X(net2669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2634 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][38] ),
    .X(net2670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2635 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][1] ),
    .X(net2671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2636 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][4] ),
    .X(net2672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2637 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ),
    .X(net2673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2638 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][35] ),
    .X(net2674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2639 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][18] ),
    .X(net2675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2640 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ),
    .X(net2676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2641 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][35] ),
    .X(net2677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2642 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ),
    .X(net2678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2643 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][14] ),
    .X(net2679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2644 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][30] ),
    .X(net2680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2645 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][7] ),
    .X(net2681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2646 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][38] ),
    .X(net2682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2647 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][36] ),
    .X(net2683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2648 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][43] ),
    .X(net2684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2649 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][7] ),
    .X(net2685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2650 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][37] ),
    .X(net2686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2651 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][15] ),
    .X(net2687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2652 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][3] ),
    .X(net2688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2653 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][17] ),
    .X(net2689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2654 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ),
    .X(net2690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2655 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][40] ),
    .X(net2691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2656 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ),
    .X(net2692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2657 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][12] ),
    .X(net2693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2658 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ),
    .X(net2694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2659 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][38] ),
    .X(net2695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2660 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][13] ),
    .X(net2696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2661 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ),
    .X(net2697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2662 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][13] ),
    .X(net2698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2663 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][19] ),
    .X(net2699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2664 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][30] ),
    .X(net2700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2665 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][0] ),
    .X(net2701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2666 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][6] ),
    .X(net2702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2667 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ),
    .X(net2703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2668 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][6] ),
    .X(net2704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2669 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][27] ),
    .X(net2705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2670 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][26] ),
    .X(net2706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2671 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][28] ),
    .X(net2707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2672 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ),
    .X(net2708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2673 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][1] ),
    .X(net2709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2674 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][21] ),
    .X(net2710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2675 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][6] ),
    .X(net2711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2676 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][42] ),
    .X(net2712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2677 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ),
    .X(net2713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2678 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][11] ),
    .X(net2714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2679 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][46] ),
    .X(net2715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2680 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][45] ),
    .X(net2716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2681 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ),
    .X(net2717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2682 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][39] ),
    .X(net2718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2683 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][0] ),
    .X(net2719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2684 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][14] ),
    .X(net2720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2685 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][1] ),
    .X(net2721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2686 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][42] ),
    .X(net2722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2687 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[1][34] ),
    .X(net2723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2688 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][34] ),
    .X(net2724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2689 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ),
    .X(net2725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2690 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ),
    .X(net2726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2691 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][3] ),
    .X(net2727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2692 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][12] ),
    .X(net2728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2693 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ),
    .X(net2729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2694 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][39] ),
    .X(net2730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2695 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][13] ),
    .X(net2731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2696 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][5] ),
    .X(net2732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2697 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][25] ),
    .X(net2733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2698 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][1] ),
    .X(net2734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2699 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ),
    .X(net2735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2700 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][30] ),
    .X(net2736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2701 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][43] ),
    .X(net2737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2702 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ),
    .X(net2738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2703 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][12] ),
    .X(net2739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2704 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][5] ),
    .X(net2740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2705 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ),
    .X(net2741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2706 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][19] ),
    .X(net2742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2707 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][32] ),
    .X(net2743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2708 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][25] ),
    .X(net2744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2709 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][41] ),
    .X(net2745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2710 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ),
    .X(net2746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2711 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][34] ),
    .X(net2747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2712 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][5] ),
    .X(net2748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2713 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][4] ),
    .X(net2749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2714 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][23] ),
    .X(net2750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2715 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][11] ),
    .X(net2751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2716 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][43] ),
    .X(net2752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2717 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][12] ),
    .X(net2753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2718 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][46] ),
    .X(net2754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2719 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][24] ),
    .X(net2755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2720 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ),
    .X(net2756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2721 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][7] ),
    .X(net2757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2722 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][32] ),
    .X(net2758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2723 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][5] ),
    .X(net2759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2724 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][17] ),
    .X(net2760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2725 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][41] ),
    .X(net2761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2726 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][34] ),
    .X(net2762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2727 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][12] ),
    .X(net2763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2728 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][5] ),
    .X(net2764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2729 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][16] ),
    .X(net2765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2730 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][20] ),
    .X(net2766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2731 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][14] ),
    .X(net2767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2732 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][7] ),
    .X(net2768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2733 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][23] ),
    .X(net2769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2734 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][29] ),
    .X(net2770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2735 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][40] ),
    .X(net2771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2736 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][3] ),
    .X(net2772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2737 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][41] ),
    .X(net2773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2738 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][29] ),
    .X(net2774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2739 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][9] ),
    .X(net2775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2740 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][8] ),
    .X(net2776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2741 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][29] ),
    .X(net2777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2742 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][33] ),
    .X(net2778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2743 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][4] ),
    .X(net2779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2744 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][2] ),
    .X(net2780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2745 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][41] ),
    .X(net2781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2746 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][37] ),
    .X(net2782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2747 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][10] ),
    .X(net2783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2748 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][4] ),
    .X(net2784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2749 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][16] ),
    .X(net2785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2750 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][26] ),
    .X(net2786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2751 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][34] ),
    .X(net2787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2752 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[0][9] ),
    .X(net2788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2753 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][9] ),
    .X(net2789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2754 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][39] ),
    .X(net2790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2755 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][0] ),
    .X(net2791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2756 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][34] ),
    .X(net2792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2757 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][14] ),
    .X(net2793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2758 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][2] ),
    .X(net2794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2759 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][29] ),
    .X(net2795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2760 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][27] ),
    .X(net2796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2761 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][42] ),
    .X(net2797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2762 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][44] ),
    .X(net2798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2763 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][33] ),
    .X(net2799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2764 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[2][10] ),
    .X(net2800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2765 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][28] ),
    .X(net2801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2766 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][10] ),
    .X(net2802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2767 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ),
    .X(net2803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2768 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][46] ),
    .X(net2804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2769 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][26] ),
    .X(net2805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2770 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][6] ),
    .X(net2806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2771 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][28] ),
    .X(net2807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2772 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][40] ),
    .X(net2808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2773 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][33] ),
    .X(net2809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2774 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][13] ),
    .X(net2810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2775 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][37] ),
    .X(net2811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2776 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ),
    .X(net2812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2777 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ),
    .X(net2813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2778 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][8] ),
    .X(net2814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2779 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][9] ),
    .X(net2815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2780 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][23] ),
    .X(net2816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2781 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][46] ),
    .X(net2817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2782 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][26] ),
    .X(net2818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2783 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][15] ),
    .X(net2819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2784 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ),
    .X(net2820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2785 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][26] ),
    .X(net2821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2786 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][13] ),
    .X(net2822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2787 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][21] ),
    .X(net2823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2788 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][19] ),
    .X(net2824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2789 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][27] ),
    .X(net2825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2790 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][21] ),
    .X(net2826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2791 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][33] ),
    .X(net2827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2792 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][14] ),
    .X(net2828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2793 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][25] ),
    .X(net2829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2794 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][32] ),
    .X(net2830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2795 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][27] ),
    .X(net2831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2796 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][41] ),
    .X(net2832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2797 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][38] ),
    .X(net2833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2798 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][2] ),
    .X(net2834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2799 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ),
    .X(net2835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2800 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][44] ),
    .X(net2836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2801 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ),
    .X(net2837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2802 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][30] ),
    .X(net2838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2803 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][43] ),
    .X(net2839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2804 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][44] ),
    .X(net2840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2805 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][36] ),
    .X(net2841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2806 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][28] ),
    .X(net2842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2807 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][31] ),
    .X(net2843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2808 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][28] ),
    .X(net2844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2809 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][23] ),
    .X(net2845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2810 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][18] ),
    .X(net2846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2811 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][13] ),
    .X(net2847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2812 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][20] ),
    .X(net2848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2813 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][38] ),
    .X(net2849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2814 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][20] ),
    .X(net2850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2815 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][41] ),
    .X(net2851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2816 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][18] ),
    .X(net2852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2817 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][24] ),
    .X(net2853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2818 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][28] ),
    .X(net2854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2819 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][34] ),
    .X(net2855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2820 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][3] ),
    .X(net2856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2821 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][35] ),
    .X(net2857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2822 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][38] ),
    .X(net2858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2823 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][15] ),
    .X(net2859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2824 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[0][7] ),
    .X(net2860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2825 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][25] ),
    .X(net2861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2826 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ),
    .X(net2862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2827 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][30] ),
    .X(net2863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2828 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][17] ),
    .X(net2864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2829 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][0] ),
    .X(net2865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2830 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[1][24] ),
    .X(net2866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2831 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][4] ),
    .X(net2867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2832 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ),
    .X(net2868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2833 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ),
    .X(net2869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2834 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][1] ),
    .X(net2870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2835 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][21] ),
    .X(net2871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2836 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][30] ),
    .X(net2872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2837 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][17] ),
    .X(net2873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2838 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][9] ),
    .X(net2874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2839 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][44] ),
    .X(net2875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2840 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[1][21] ),
    .X(net2876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2841 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][41] ),
    .X(net2877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2842 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ),
    .X(net2878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2843 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][4] ),
    .X(net2879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2844 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][0] ),
    .X(net2880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2845 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][3] ),
    .X(net2881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2846 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][19] ),
    .X(net2882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2847 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][9] ),
    .X(net2883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2848 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][7] ),
    .X(net2884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2849 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][46] ),
    .X(net2885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2850 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][28] ),
    .X(net2886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2851 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][12] ),
    .X(net2887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2852 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ),
    .X(net2888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2853 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][21] ),
    .X(net2889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2854 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][17] ),
    .X(net2890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2855 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][40] ),
    .X(net2891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2856 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][9] ),
    .X(net2892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2857 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][32] ),
    .X(net2893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2858 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][0] ),
    .X(net2894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2859 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ),
    .X(net2895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2860 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][3] ),
    .X(net2896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2861 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][35] ),
    .X(net2897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2862 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][3] ),
    .X(net2898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2863 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][22] ),
    .X(net2899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2864 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][29] ),
    .X(net2900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2865 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.ram[1][25] ),
    .X(net2901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2866 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ),
    .X(net2902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2867 (.A(\c.genblk1.genblk1.subs.sw.up.x.o[2] ),
    .X(net2903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2868 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .X(net2904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2869 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.ram[0][13] ),
    .X(net2905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2870 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][8] ),
    .X(net2906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2871 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][8] ),
    .X(net2907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2872 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][11] ),
    .X(net2908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2873 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[1][20] ),
    .X(net2909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2874 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][15] ),
    .X(net2910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2875 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[0][25] ),
    .X(net2911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2876 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][42] ),
    .X(net2912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2877 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][39] ),
    .X(net2913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2878 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][12] ),
    .X(net2914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2879 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][22] ),
    .X(net2915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2880 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[0][29] ),
    .X(net2916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2881 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[2][24] ),
    .X(net2917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2882 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ),
    .X(net2918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2883 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][46] ),
    .X(net2919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2884 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[0][22] ),
    .X(net2920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2885 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][2] ),
    .X(net2921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2886 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ),
    .X(net2922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2887 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][15] ),
    .X(net2923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2888 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][46] ),
    .X(net2924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2889 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ),
    .X(net2925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2890 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][20] ),
    .X(net2926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2891 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][38] ),
    .X(net2927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2892 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][40] ),
    .X(net2928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2893 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.ram[2][30] ),
    .X(net2929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2894 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][14] ),
    .X(net2930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2895 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][2] ),
    .X(net2931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2896 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][40] ),
    .X(net2932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2897 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][37] ),
    .X(net2933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2898 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][20] ),
    .X(net2934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2899 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.ram[1][32] ),
    .X(net2935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2900 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][26] ),
    .X(net2936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2901 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][22] ),
    .X(net2937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2902 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][0] ),
    .X(net2938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2903 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ),
    .X(net2939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2904 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[0][26] ),
    .X(net2940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2905 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .X(net2941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2906 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][22] ),
    .X(net2942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2907 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][36] ),
    .X(net2943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2908 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][21] ),
    .X(net2944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2909 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][14] ),
    .X(net2945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2910 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .X(net2946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2911 (.A(\c.genblk1.genblk1.subs.sw.up.x.o[1] ),
    .X(net2947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2912 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .X(net2948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2913 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[2][5] ),
    .X(net2949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2914 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.ram[2][28] ),
    .X(net2950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2915 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .X(net2951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2916 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .X(net2952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2917 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][31] ),
    .X(net2953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2918 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .X(net2954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2919 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .X(net2955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2920 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .X(net2956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2921 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .X(net2957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2922 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .X(net2958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2923 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .X(net2959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2924 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .X(net2960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2925 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .X(net2961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2926 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .X(net2962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2927 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .X(net2963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2928 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .X(net2964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2929 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .X(net2965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2930 (.A(\c.cfg_i_q[2] ),
    .X(net2966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2931 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .X(net2967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2932 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .X(net2968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2933 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .X(net2969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2934 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .X(net2970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2935 (.A(\c.genblk1.genblk1.subs.sw.up.x.o[0] ),
    .X(net2971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2936 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .X(net2972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2937 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .X(net2973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2938 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .X(net2974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2939 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .X(net2975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2940 (.A(\c.genblk1.genblk1.subs.sw.up.x.o[6] ),
    .X(net2976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2941 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .X(net2977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2942 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .X(net2978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2943 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .X(net2979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2944 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ),
    .X(net2980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2945 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .X(net2981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2946 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .X(net2982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2947 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .X(net2983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2948 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .X(net2984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2949 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .X(net2985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2950 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .X(net2986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2951 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .X(net2987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2952 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .X(net2988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2953 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .X(net2989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2954 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .X(net2990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2955 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .X(net2991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2956 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .X(net2992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2957 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .X(net2993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2958 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .X(net2994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2959 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .X(net2995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2960 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .X(net2996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2961 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .X(net2997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2962 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .X(net2998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2963 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .X(net2999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2964 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ),
    .X(net3000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2965 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .X(net3001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2966 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .X(net3002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2967 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .X(net3003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2968 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .X(net3004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2969 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .X(net3005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2970 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .X(net3006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2971 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .X(net3007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2972 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .X(net3008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2973 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .X(net3009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2974 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .X(net3010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2975 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .X(net3011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2976 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .X(net3012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2977 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .X(net3013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2978 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .X(net3014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2979 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .X(net3015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2980 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .X(net3016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2981 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .X(net3017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2982 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .X(net3018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2983 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .X(net3019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2984 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .X(net3020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2985 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .X(net3021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2986 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .X(net3022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2987 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .X(net3023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2988 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[10] ),
    .X(net3024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2989 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .X(net3025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2990 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .X(net3026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2991 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .X(net3027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2992 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .X(net3028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2993 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .X(net3029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2994 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .X(net3030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2995 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .X(net3031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2996 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .X(net3032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2997 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .X(net3033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2998 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .X(net3034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2999 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .X(net3035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3000 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .X(net3036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3001 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .X(net3037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3002 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .X(net3038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3003 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .X(net3039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3004 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .X(net3040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3005 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[4] ),
    .X(net3041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3006 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .X(net3042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3007 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .X(net3043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3008 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .X(net3044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3009 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[5] ),
    .X(net3045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3010 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[9] ),
    .X(net3046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3011 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .X(net3047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3012 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .X(net3048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3013 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .X(net3049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3014 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .X(net3050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3015 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[2] ),
    .X(net3051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3016 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .X(net3052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3017 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .X(net3053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3018 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .X(net3054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3019 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .X(net3055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3020 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .X(net3056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3021 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .X(net3057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3022 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .X(net3058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3023 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[1] ),
    .X(net3059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3024 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .X(net3060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3025 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .X(net3061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3026 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .X(net3062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3027 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .X(net3063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3028 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .X(net3064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3029 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .X(net3065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3030 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[10] ),
    .X(net3066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3031 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .X(net3067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3032 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .X(net3068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3033 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .X(net3069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3034 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[1] ),
    .X(net3070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3035 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[5] ),
    .X(net3071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3036 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .X(net3072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3037 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .X(net3073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3038 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[1] ),
    .X(net3074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3039 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ),
    .X(net3075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3040 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[5] ),
    .X(net3076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3041 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[10] ),
    .X(net3077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3042 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[9] ),
    .X(net3078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3043 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[6] ),
    .X(net3079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3044 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .X(net3080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3045 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .X(net3081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3046 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .X(net3082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3047 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[2] ),
    .X(net3083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3048 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[2] ),
    .X(net3084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3049 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .X(net3085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3050 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .X(net3086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3051 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .X(net3087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3052 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .X(net3088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3053 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .X(net3089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3054 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[6] ),
    .X(net3090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3055 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[2][28] ),
    .X(net3091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3056 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[6] ),
    .X(net3092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3057 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .X(net3093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3058 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .X(net3094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3059 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .X(net3095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3060 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[5] ),
    .X(net3096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3061 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[4] ),
    .X(net3097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3062 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[9] ),
    .X(net3098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3063 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[1] ),
    .X(net3099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3064 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.ram[1][29] ),
    .X(net3100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3065 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .X(net3101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3066 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .X(net3102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3067 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ),
    .X(net3103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3068 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .X(net3104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3069 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .X(net3105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3070 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .X(net3106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3071 (.A(\c.genblk1.genblk1.subs.sw.up.x.o[5] ),
    .X(net3107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3072 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.ram[0][32] ),
    .X(net3108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3073 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[9] ),
    .X(net3109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3074 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .X(net3110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3075 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[14] ),
    .X(net3111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3076 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[10] ),
    .X(net3112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3077 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .X(net3113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3078 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][17] ),
    .X(net3114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3079 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ),
    .X(net3115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3080 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .X(net3116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3081 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][16] ),
    .X(net3117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3082 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[14] ),
    .X(net3118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3083 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ),
    .X(net3119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3084 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[13] ),
    .X(net3120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3085 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ),
    .X(net3121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3086 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[13] ),
    .X(net3122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3087 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .X(net3123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3088 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ),
    .X(net3124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3089 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[14] ),
    .X(net3125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3090 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .X(net3126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3091 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[14] ),
    .X(net3127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3092 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ),
    .X(net3128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3093 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ),
    .X(net3129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3094 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[13] ),
    .X(net3130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3095 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .X(net3131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3096 (.A(_03421_),
    .X(net3132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3097 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fds ),
    .X(net3133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3098 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[13] ),
    .X(net3134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3099 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .X(net3135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3100 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ),
    .X(net3136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3101 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[8] ),
    .X(net3137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3102 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .X(net3138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3103 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ),
    .X(net3139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3104 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ),
    .X(net3140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3105 (.A(_01148_),
    .X(net3141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3106 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[22] ),
    .X(net3142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3107 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ),
    .X(net3143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3108 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ),
    .X(net3144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3109 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ),
    .X(net3145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3110 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fds ),
    .X(net3146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3111 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ),
    .X(net3147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3112 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ),
    .X(net3148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3113 (.A(_01233_),
    .X(net3149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3114 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ),
    .X(net3150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3115 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ),
    .X(net3151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3116 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ),
    .X(net3152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3117 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .X(net3153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3118 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ),
    .X(net3154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3119 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .X(net3155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3120 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ),
    .X(net3156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3121 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ),
    .X(net3157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3122 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .X(net3158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3123 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ),
    .X(net3159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3124 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ),
    .X(net3160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3125 (.A(_02523_),
    .X(net3161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3126 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ),
    .X(net3162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3127 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .X(net3163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3128 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ),
    .X(net3164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3129 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ),
    .X(net3165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3130 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .X(net3166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3131 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ),
    .X(net3167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3132 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[14] ),
    .X(net3168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3133 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[27] ),
    .X(net3169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3134 (.A(\c.genblk1.genblk1.subs.sw.up.x.o_[6] ),
    .X(net3170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3135 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ),
    .X(net3171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3136 (.A(_00795_),
    .X(net3172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3137 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ),
    .X(net3173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3138 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ),
    .X(net3174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3139 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .X(net3175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3140 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ),
    .X(net3176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3141 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ),
    .X(net3177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3142 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[6] ),
    .X(net3178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3143 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ),
    .X(net3179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3144 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[0] ),
    .X(net3180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3145 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .X(net3181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3146 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ),
    .X(net3182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3147 (.A(_00142_),
    .X(net3183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3148 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[0] ),
    .X(net3184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3149 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[15] ),
    .X(net3185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3150 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .X(net3186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3151 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fds ),
    .X(net3187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3152 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ),
    .X(net3188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3153 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ),
    .X(net3189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3154 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[0] ),
    .X(net3190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3155 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[19] ),
    .X(net3191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3156 (.A(\c.genblk1.genblk1.subs.sw.up.x.o_[4] ),
    .X(net3192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3157 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ),
    .X(net3193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3158 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .X(net3194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3159 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ),
    .X(net3195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3160 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .X(net3196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3161 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ),
    .X(net3197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3162 (.A(_02747_),
    .X(net3198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3163 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[0] ),
    .X(net3199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3164 (.A(_04582_),
    .X(net3200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3165 (.A(_00046_),
    .X(net3201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3166 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ),
    .X(net3202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3167 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .X(net3203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3168 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ),
    .X(net3204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3169 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .X(net3205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3170 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ),
    .X(net3206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3171 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ),
    .X(net3207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3172 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ),
    .X(net3208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3173 (.A(_00097_),
    .X(net3209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3174 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .X(net3210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3175 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .X(net3211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3176 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .X(net3212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3177 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ),
    .X(net3213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3178 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ),
    .X(net3214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3179 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[7] ),
    .X(net3215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3180 (.A(\c.genblk1.genblk1.subs.sw.up.x.o_[1] ),
    .X(net3216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3181 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(net3217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3182 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.fds ),
    .X(net3218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3183 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ),
    .X(net3219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3184 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ),
    .X(net3220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3185 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ),
    .X(net3221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3186 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ),
    .X(net3222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3187 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ),
    .X(net3223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3188 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ),
    .X(net3224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3189 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[3] ),
    .X(net3225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3190 (.A(\c.genblk1.genblk1.subs.sw.up.x.o_[0] ),
    .X(net3226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3191 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .X(net3227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3192 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fds ),
    .X(net3228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3193 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ),
    .X(net3229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3194 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ),
    .X(net3230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3195 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.fds ),
    .X(net3231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3196 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ),
    .X(net3232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3197 (.A(_02328_),
    .X(net3233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3198 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fds ),
    .X(net3234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3199 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[45] ),
    .X(net3235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3200 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .X(net3236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3201 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ),
    .X(net3237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3202 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ),
    .X(net3238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3203 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .X(net3239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3204 (.A(_04595_),
    .X(net3240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3205 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .X(net3241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3206 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fds ),
    .X(net3242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3207 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .X(net3243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3208 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ),
    .X(net3244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3209 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[12] ),
    .X(net3245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3210 (.A(_03858_),
    .X(net3246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3211 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[1] ),
    .X(net3247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3212 (.A(_04553_),
    .X(net3248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3213 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(net3249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3214 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .X(net3250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3215 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(net3251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3216 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .X(net3252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3217 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .X(net3253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3218 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ),
    .X(net3254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3219 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[0] ),
    .X(net3255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3220 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[24] ),
    .X(net3256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3221 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[0] ),
    .X(net3257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3222 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ),
    .X(net3258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3223 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fde ),
    .X(net3259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3224 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.fde ),
    .X(net3260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3225 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ),
    .X(net3261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3226 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ),
    .X(net3262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3227 (.A(_01870_),
    .X(net3263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3228 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(net3264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3229 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(net3265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3230 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ),
    .X(net3266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3231 (.A(_04681_),
    .X(net3267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3232 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .X(net3268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3233 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(net3269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3234 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(net3270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3235 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .X(net3271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3236 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[44] ),
    .X(net3272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3237 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ),
    .X(net3273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3238 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ),
    .X(net3274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3239 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .X(net3275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3240 (.A(_00165_),
    .X(net3276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3241 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(net3277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3242 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .X(net3278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3243 (.A(_04652_),
    .X(net3279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3244 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(net3280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3245 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ),
    .X(net3281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3246 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[22] ),
    .X(net3282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3247 (.A(_04264_),
    .X(net3283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3248 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[4] ),
    .X(net3284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3249 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ),
    .X(net3285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3250 (.A(_01314_),
    .X(net3286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3251 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[9] ),
    .X(net3287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3252 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[1] ),
    .X(net3288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3253 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .X(net3289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3254 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .X(net3290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3255 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[1] ),
    .X(net3291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3256 (.A(_02529_),
    .X(net3292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3257 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ),
    .X(net3293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3258 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[0] ),
    .X(net3294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3259 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .X(net3295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3260 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ),
    .X(net3296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3261 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .X(net3297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3262 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .X(net3298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3263 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ),
    .X(net3299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3264 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ),
    .X(net3300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3265 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ),
    .X(net3301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3266 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ),
    .X(net3302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3267 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .X(net3303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3268 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[1] ),
    .X(net3304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3269 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .X(net3305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3270 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.sr.ram_in[46] ),
    .X(net3306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3271 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[39] ),
    .X(net3307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3272 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[7] ),
    .X(net3308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3273 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[29] ),
    .X(net3309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3274 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ),
    .X(net3310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3275 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .X(net3311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3276 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ),
    .X(net3312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3277 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .X(net3313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3278 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fde ),
    .X(net3314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3279 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ),
    .X(net3315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3280 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ),
    .X(net3316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3281 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[34] ),
    .X(net3317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3282 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ),
    .X(net3318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3283 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ),
    .X(net3319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3284 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ),
    .X(net3320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3285 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ),
    .X(net3321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3286 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.fd ),
    .X(net3322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3287 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .X(net3323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3288 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ),
    .X(net3324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3289 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ),
    .X(net3325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3290 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ),
    .X(net3326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3291 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ),
    .X(net3327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3292 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ),
    .X(net3328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3293 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ),
    .X(net3329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3294 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(net3330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3295 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ),
    .X(net3331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3296 (.A(_02532_),
    .X(net3332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3297 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ),
    .X(net3333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3298 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ),
    .X(net3334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3299 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[1] ),
    .X(net3335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3300 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ),
    .X(net3336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3301 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ),
    .X(net3337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3302 (.A(_03328_),
    .X(net3338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3303 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ),
    .X(net3339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3304 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.fd ),
    .X(net3340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3305 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[13] ),
    .X(net3341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3306 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ),
    .X(net3342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3307 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ),
    .X(net3343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3308 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ),
    .X(net3344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3309 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ),
    .X(net3345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3310 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ),
    .X(net3346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3311 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ),
    .X(net3347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3312 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .X(net3348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3313 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ),
    .X(net3349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3314 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ),
    .X(net3350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3315 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ),
    .X(net3351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3316 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ),
    .X(net3352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3317 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ),
    .X(net3353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3318 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[15] ),
    .X(net3354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3319 (.A(\c.genblk1.genblk1.subs.sw.up.x.o_[3] ),
    .X(net3355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3320 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ),
    .X(net3356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3321 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ),
    .X(net3357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3322 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ),
    .X(net3358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3323 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ),
    .X(net3359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3324 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ),
    .X(net3360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3325 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ),
    .X(net3361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3326 (.A(_02754_),
    .X(net3362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3327 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ),
    .X(net3363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3328 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ),
    .X(net3364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3329 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ),
    .X(net3365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3330 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ),
    .X(net3366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3331 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[1] ),
    .X(net3367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3332 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ),
    .X(net3368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3333 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ),
    .X(net3369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3334 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ),
    .X(net3370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3335 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .X(net3371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3336 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .X(net3372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3337 (.A(_03097_),
    .X(net3373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3338 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .X(net3374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3339 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .X(net3375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3340 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .X(net3376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3341 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[1] ),
    .X(net3377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3342 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[1] ),
    .X(net3378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3343 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.fde ),
    .X(net3379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3344 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ),
    .X(net3380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3345 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ),
    .X(net3381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3346 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .X(net3382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3347 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ),
    .X(net3383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3348 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ),
    .X(net3384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3349 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ),
    .X(net3385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3350 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ),
    .X(net3386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3351 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ),
    .X(net3387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3352 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[11] ),
    .X(net3388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3353 (.A(\c.genblk1.genblk1.subs.sw.up.x.o_[2] ),
    .X(net3389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3354 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[24] ),
    .X(net3390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3355 (.A(_03581_),
    .X(net3391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3356 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[4] ),
    .X(net3392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3357 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ),
    .X(net3393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3358 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ),
    .X(net3394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3359 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[14] ),
    .X(net3395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3360 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ),
    .X(net3396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3361 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ),
    .X(net3397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3362 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ),
    .X(net3398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3363 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ),
    .X(net3399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3364 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .X(net3400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3365 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ),
    .X(net3401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3366 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ),
    .X(net3402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3367 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ),
    .X(net3403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3368 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ),
    .X(net3404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3369 (.A(_01877_),
    .X(net3405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3370 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(net3406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3371 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ),
    .X(net3407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3372 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.fd ),
    .X(net3408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3373 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ),
    .X(net3409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3374 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ),
    .X(net3410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3375 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ),
    .X(net3411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3376 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ),
    .X(net3412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3377 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ),
    .X(net3413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3378 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ),
    .X(net3414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3379 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[4] ),
    .X(net3415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3380 (.A(_03737_),
    .X(net3416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3381 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[0] ),
    .X(net3417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3382 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[10] ),
    .X(net3418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3383 (.A(_01414_),
    .X(net3419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3384 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ),
    .X(net3420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3385 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ),
    .X(net3421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3386 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[8] ),
    .X(net3422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3387 (.A(_04092_),
    .X(net3423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3388 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[1] ),
    .X(net3424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3389 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[4] ),
    .X(net3425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3390 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(net3426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3391 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ),
    .X(net3427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3392 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ),
    .X(net3428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3393 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ),
    .X(net3429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3394 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ),
    .X(net3430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3395 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .X(net3431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3396 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ),
    .X(net3432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3397 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[19] ),
    .X(net3433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3398 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[5] ),
    .X(net3434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3399 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ),
    .X(net3435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3400 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ),
    .X(net3436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3401 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ),
    .X(net3437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3402 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ),
    .X(net3438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3403 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ),
    .X(net3439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3404 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ),
    .X(net3440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3405 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ),
    .X(net3441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3406 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ),
    .X(net3442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3407 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .X(net3443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3408 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ),
    .X(net3444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3409 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ),
    .X(net3445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3410 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .X(net3446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3411 (.A(_00159_),
    .X(net3447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3412 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ),
    .X(net3448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3413 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ),
    .X(net3449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3414 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ),
    .X(net3450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3415 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ),
    .X(net3451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3416 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .X(net3452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3417 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ),
    .X(net3453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3418 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ),
    .X(net3454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3419 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ),
    .X(net3455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3420 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ),
    .X(net3456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3421 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ),
    .X(net3457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3422 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ),
    .X(net3458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3423 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ),
    .X(net3459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3424 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ),
    .X(net3460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3425 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ),
    .X(net3461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3426 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ),
    .X(net3462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3427 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .X(net3463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3428 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ),
    .X(net3464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3429 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ),
    .X(net3465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3430 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ),
    .X(net3466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3431 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ),
    .X(net3467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3432 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ),
    .X(net3468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3433 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ),
    .X(net3469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3434 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[0] ),
    .X(net3470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3435 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(net3471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3436 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[12] ),
    .X(net3472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3437 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .X(net3473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3438 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[14] ),
    .X(net3474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3439 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .X(net3475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3440 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ),
    .X(net3476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3441 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ),
    .X(net3477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3442 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ),
    .X(net3478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3443 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ),
    .X(net3479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3444 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ),
    .X(net3480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3445 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ),
    .X(net3481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3446 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(net3482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3447 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ),
    .X(net3483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3448 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ),
    .X(net3484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3449 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ),
    .X(net3485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3450 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ),
    .X(net3486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3451 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[12] ),
    .X(net3487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3452 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[9] ),
    .X(net3488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3453 (.A(_03696_),
    .X(net3489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3454 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[1] ),
    .X(net3490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3455 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ),
    .X(net3491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3456 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(net3492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3457 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .X(net3493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3458 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[29] ),
    .X(net3494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3459 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[5] ),
    .X(net3495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3460 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ),
    .X(net3496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3461 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ),
    .X(net3497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3462 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ),
    .X(net3498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3463 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ),
    .X(net3499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3464 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[1] ),
    .X(net3500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3465 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ),
    .X(net3501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3466 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .X(net3502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3467 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ),
    .X(net3503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3468 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[39] ),
    .X(net3504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3469 (.A(_04000_),
    .X(net3505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3470 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[7] ),
    .X(net3506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3471 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[12] ),
    .X(net3507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3472 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ),
    .X(net3508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3473 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ),
    .X(net3509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3474 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[5] ),
    .X(net3510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3475 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[2] ),
    .X(net3511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3476 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[3] ),
    .X(net3512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3477 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ),
    .X(net3513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3478 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .X(net3514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3479 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[5] ),
    .X(net3515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3480 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ),
    .X(net3516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3481 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .X(net3517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3482 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ),
    .X(net3518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3483 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ),
    .X(net3519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3484 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ),
    .X(net3520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3485 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ),
    .X(net3521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3486 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ),
    .X(net3522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3487 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ),
    .X(net3523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3488 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ),
    .X(net3524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3489 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ),
    .X(net3525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3490 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[14] ),
    .X(net3526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3491 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ),
    .X(net3527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3492 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[3] ),
    .X(net3528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3493 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[1] ),
    .X(net3529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3494 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[14] ),
    .X(net3530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3495 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ),
    .X(net3531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3496 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ),
    .X(net3532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3497 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .X(net3533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3498 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[4] ),
    .X(net3534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3499 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .X(net3535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3500 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[6] ),
    .X(net3536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3501 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[2] ),
    .X(net3537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3502 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[37] ),
    .X(net3538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3503 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .X(net3539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3504 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ),
    .X(net3540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3505 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ),
    .X(net3541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3506 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ),
    .X(net3542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3507 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ),
    .X(net3543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3508 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ),
    .X(net3544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3509 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ),
    .X(net3545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3510 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[12] ),
    .X(net3546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3511 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ),
    .X(net3547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3512 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .X(net3548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3513 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ),
    .X(net3549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3514 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .X(net3550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3515 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ),
    .X(net3551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3516 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .X(net3552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3517 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ),
    .X(net3553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3518 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[4] ),
    .X(net3554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3519 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ),
    .X(net3555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3520 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ),
    .X(net3556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3521 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ),
    .X(net3557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3522 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ),
    .X(net3558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3523 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ),
    .X(net3559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3524 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ),
    .X(net3560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3525 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[14] ),
    .X(net3561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3526 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ),
    .X(net3562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3527 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ),
    .X(net3563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3528 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ),
    .X(net3564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3529 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[5] ),
    .X(net3565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3530 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[4] ),
    .X(net3566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3531 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[15] ),
    .X(net3567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3532 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ),
    .X(net3568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3533 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ),
    .X(net3569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3534 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ),
    .X(net3570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3535 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ),
    .X(net3571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3536 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ),
    .X(net3572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3537 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[5] ),
    .X(net3573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3538 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[4] ),
    .X(net3574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3539 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[29] ),
    .X(net3575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3540 (.A(_03814_),
    .X(net3576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3541 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[5] ),
    .X(net3577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3542 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[6] ),
    .X(net3578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3543 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ),
    .X(net3579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3544 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ),
    .X(net3580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3545 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .X(net3581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3546 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[13] ),
    .X(net3582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3547 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .X(net3583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3548 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(net3584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3549 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ),
    .X(net3585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3550 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[5] ),
    .X(net3586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3551 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[3] ),
    .X(net3587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3552 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ),
    .X(net3588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3553 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[7] ),
    .X(net3589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3554 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ),
    .X(net3590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3555 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[13] ),
    .X(net3591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3556 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .X(net3592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3557 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ),
    .X(net3593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3558 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[14] ),
    .X(net3594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3559 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .X(net3595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3560 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .X(net3596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3561 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .X(net3597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3562 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[29] ),
    .X(net3598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3563 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(net3599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3564 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .X(net3600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3565 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ),
    .X(net3601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3566 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ),
    .X(net3602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3567 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ),
    .X(net3603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3568 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ),
    .X(net3604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3569 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ),
    .X(net3605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3570 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ),
    .X(net3606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3571 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[10] ),
    .X(net3607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3572 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .X(net3608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3573 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[7] ),
    .X(net3609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3574 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(net3610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3575 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ),
    .X(net3611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3576 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[15] ),
    .X(net3612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3577 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[0] ),
    .X(net3613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3578 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ),
    .X(net3614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3579 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[15] ),
    .X(net3615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3580 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ),
    .X(net3616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3581 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ),
    .X(net3617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3582 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[9] ),
    .X(net3618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3583 (.A(_03899_),
    .X(net3619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3584 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[1] ),
    .X(net3620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3585 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .X(net3621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3586 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[13] ),
    .X(net3622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3587 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[5] ),
    .X(net3623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3588 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ),
    .X(net3624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3589 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[5] ),
    .X(net3625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3590 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ),
    .X(net3626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3591 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ),
    .X(net3627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3592 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ),
    .X(net3628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3593 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .X(net3629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3594 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ),
    .X(net3630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3595 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[39] ),
    .X(net3631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3596 (.A(_03483_),
    .X(net3632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3597 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[7] ),
    .X(net3633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3598 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ),
    .X(net3634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3599 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .X(net3635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3600 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(net3636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3601 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .X(net3637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3602 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .X(net3638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3603 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[7] ),
    .X(net3639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3604 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ),
    .X(net3640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3605 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ),
    .X(net3641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3606 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[9] ),
    .X(net3642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3607 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .X(net3643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3608 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .X(net3644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3609 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[7] ),
    .X(net3645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3610 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[31] ),
    .X(net3646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3611 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .X(net3647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3612 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ),
    .X(net3648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3613 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(net3649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3614 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[30] ),
    .X(net3650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3615 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ),
    .X(net3651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3616 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[5] ),
    .X(net3652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3617 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .X(net3653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3618 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ),
    .X(net3654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3619 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[10] ),
    .X(net3655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3620 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ),
    .X(net3656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3621 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.fd ),
    .X(net3657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3622 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ),
    .X(net3658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3623 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ),
    .X(net3659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3624 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(net3660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3625 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[5] ),
    .X(net3661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3626 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[15] ),
    .X(net3662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3627 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[14] ),
    .X(net3663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3628 (.A(_03658_),
    .X(net3664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3629 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.o_[2] ),
    .X(net3665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3630 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[1] ),
    .X(net3666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3631 (.A(\c.genblk1.genblk1.subs.c0.cfg_i_q[2] ),
    .X(net3667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3632 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ),
    .X(net3668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3633 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .X(net3669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3634 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(net3670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3635 (.A(_00145_),
    .X(net3671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3636 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[2] ),
    .X(net3672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3637 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ),
    .X(net3673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3638 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .X(net3674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3639 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ),
    .X(net3675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3640 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[1] ),
    .X(net3676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3641 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[19] ),
    .X(net3677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3642 (.A(_03842_),
    .X(net3678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3643 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[3] ),
    .X(net3679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3644 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[4] ),
    .X(net3680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3645 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[7] ),
    .X(net3681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3646 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ),
    .X(net3682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3647 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[13] ),
    .X(net3683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3648 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[10] ),
    .X(net3684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3649 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(net3685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3650 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ),
    .X(net3686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3651 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .X(net3687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3652 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[4] ),
    .X(net3688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3653 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[0] ),
    .X(net3689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3654 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ),
    .X(net3690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3655 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[7] ),
    .X(net3691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3656 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .X(net3692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3657 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .X(net3693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3658 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ),
    .X(net3694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3659 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .X(net3695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3660 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[4] ),
    .X(net3696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3661 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .X(net3697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3662 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .X(net3698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3663 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ),
    .X(net3699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3664 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[24] ),
    .X(net3700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3665 (.A(_03832_),
    .X(net3701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3666 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[4] ),
    .X(net3702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3667 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ),
    .X(net3703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3668 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ),
    .X(net3704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3669 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[1] ),
    .X(net3705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3670 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[1] ),
    .X(net3706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3671 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[5] ),
    .X(net3707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3672 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .X(net3708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3673 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ),
    .X(net3709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3674 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ),
    .X(net3710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3675 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ),
    .X(net3711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3676 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .X(net3712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3677 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[2] ),
    .X(net3713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3678 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .X(net3714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3679 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[24] ),
    .X(net3715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3680 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ),
    .X(net3716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3681 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ),
    .X(net3717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3682 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[10] ),
    .X(net3718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3683 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ),
    .X(net3719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3684 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[5] ),
    .X(net3720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3685 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .X(net3721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3686 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .X(net3722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3687 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ),
    .X(net3723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3688 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[34] ),
    .X(net3724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3689 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[19] ),
    .X(net3725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3690 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[5] ),
    .X(net3726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3691 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ),
    .X(net3727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3692 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[5] ),
    .X(net3728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3693 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ),
    .X(net3729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3694 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .X(net3730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3695 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ),
    .X(net3731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3696 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ),
    .X(net3732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3697 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(net3733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3698 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .X(net3734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3699 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .X(net3735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3700 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ),
    .X(net3736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3701 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[0] ),
    .X(net3737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3702 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[28] ),
    .X(net3738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3703 (.A(_04250_),
    .X(net3739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3704 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[5] ),
    .X(net3740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3705 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[10] ),
    .X(net3741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3706 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .X(net3742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3707 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[4] ),
    .X(net3743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3708 (.A(_04124_),
    .X(net3744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3709 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[0] ),
    .X(net3745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3710 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[2] ),
    .X(net3746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3711 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[10] ),
    .X(net3747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3712 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[2] ),
    .X(net3748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3713 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[3] ),
    .X(net3749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3714 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[2] ),
    .X(net3750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3715 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[7] ),
    .X(net3751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3716 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .X(net3752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3717 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[11] ),
    .X(net3753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3718 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[11] ),
    .X(net3754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3719 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[6] ),
    .X(net3755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3720 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .X(net3756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3721 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[2] ),
    .X(net3757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3722 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .X(net3758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3723 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .X(net3759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3724 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[7] ),
    .X(net3760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3725 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[4] ),
    .X(net3761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3726 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ),
    .X(net3762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3727 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .X(net3763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3728 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[34] ),
    .X(net3764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3729 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[2] ),
    .X(net3765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3730 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ),
    .X(net3766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3731 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[4] ),
    .X(net3767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3732 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ),
    .X(net3768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3733 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ),
    .X(net3769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3734 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .X(net3770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3735 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[1] ),
    .X(net3771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3736 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ),
    .X(net3772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3737 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ),
    .X(net3773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3738 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[6] ),
    .X(net3774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3739 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .X(net3775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3740 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .X(net3776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3741 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[5] ),
    .X(net3777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3742 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .X(net3778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3743 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(net3779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3744 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[8] ),
    .X(net3780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3745 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ),
    .X(net3781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3746 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .X(net3782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3747 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .X(net3783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3748 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .X(net3784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3749 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[8] ),
    .X(net3785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3750 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[3] ),
    .X(net3786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3751 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[23] ),
    .X(net3787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3752 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[32] ),
    .X(net3788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3753 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[9] ),
    .X(net3789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3754 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(net3790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3755 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ),
    .X(net3791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3756 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[7] ),
    .X(net3792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3757 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ),
    .X(net3793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3758 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(net3794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3759 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.seg[1] ),
    .X(net3795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3760 (.A(_00048_),
    .X(net3796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3761 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(net3797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3762 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .X(net3798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3763 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .X(net3799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3764 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(net3800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3765 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(net3801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3766 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .X(net3802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3767 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[4] ),
    .X(net3803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3768 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ),
    .X(net3804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3769 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[0] ),
    .X(net3805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3770 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ),
    .X(net3806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3771 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .X(net3807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3772 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ),
    .X(net3808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3773 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .X(net3809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3774 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ),
    .X(net3810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3775 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[38] ),
    .X(net3811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3776 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[11] ),
    .X(net3812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3777 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .X(net3813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3778 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[6] ),
    .X(net3814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3779 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[8] ),
    .X(net3815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3780 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[10] ),
    .X(net3816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3781 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(net3817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3782 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[37] ),
    .X(net3818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3783 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .X(net3819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3784 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_ce ),
    .X(net3820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3785 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[1] ),
    .X(net3821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3786 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[14] ),
    .X(net3822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3787 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[3] ),
    .X(net3823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3788 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[2] ),
    .X(net3824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3789 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .X(net3825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3790 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[33] ),
    .X(net3826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3791 (.A(_04234_),
    .X(net3827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3792 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[6] ),
    .X(net3828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3793 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .X(net3829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3794 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .X(net3830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3795 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[4] ),
    .X(net3831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3796 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[4] ),
    .X(net3832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3797 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ),
    .X(net3833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3798 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(net3834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3799 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ),
    .X(net3835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3800 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(net3836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3801 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[3] ),
    .X(net3837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3802 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[4] ),
    .X(net3838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3803 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .X(net3839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3804 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .X(net3840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3805 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ),
    .X(net3841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3806 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[37] ),
    .X(net3842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3807 (.A(_03766_),
    .X(net3843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3808 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.o_[7] ),
    .X(net3844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3809 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ),
    .X(net3845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3810 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(net3846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3811 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[11] ),
    .X(net3847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3812 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .X(net3848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3813 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ),
    .X(net3849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3814 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.o[8] ),
    .X(net3850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3815 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .X(net3851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3816 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .X(net3852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3817 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .X(net3853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3818 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .X(net3854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3819 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .X(net3855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3820 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[10] ),
    .X(net3856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3821 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[1] ),
    .X(net3857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3822 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[14] ),
    .X(net3858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3823 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[9] ),
    .X(net3859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3824 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(net3860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3825 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(net3861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3826 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(net3862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3827 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(net3863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3828 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(net3864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3829 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .X(net3865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3830 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[11] ),
    .X(net3866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3831 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(net3867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3832 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .X(net3868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3833 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(net3869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3834 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .X(net3870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3835 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(net3871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3836 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[2] ),
    .X(net3872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3837 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .X(net3873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3838 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[7] ),
    .X(net3874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3839 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .X(net3875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3840 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[7] ),
    .X(net3876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3841 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[4] ),
    .X(net3877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3842 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(net3878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3843 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.luts.o[8] ),
    .X(net3879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3844 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[1] ),
    .X(net3880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3845 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(net3881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3846 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[12] ),
    .X(net3882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3847 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .X(net3883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3848 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ff_rst ),
    .X(net3884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3849 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(net3885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3850 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(net3886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3851 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[5] ),
    .X(net3887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3852 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(net3888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3853 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(net3889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3854 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[19] ),
    .X(net3890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3855 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[3] ),
    .X(net3891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3856 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[2] ),
    .X(net3892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3857 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .X(net3893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3858 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(net3894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3859 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[9] ),
    .X(net3895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3860 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[12] ),
    .X(net3896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3861 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(net3897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3862 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(net3898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3863 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ),
    .X(net3899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3864 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.seg[1] ),
    .X(net3900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3865 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[14] ),
    .X(net3901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3866 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[2] ),
    .X(net3902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3867 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(net3903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3868 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .X(net3904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3869 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[10] ),
    .X(net3905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3870 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(net3906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3871 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[2] ),
    .X(net3907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3872 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(net3908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3873 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[4] ),
    .X(net3909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3874 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[6] ),
    .X(net3910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3875 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(net3911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3876 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(net3912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3877 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .X(net3913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3878 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ),
    .X(net3914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3879 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[18] ),
    .X(net3915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3880 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[9] ),
    .X(net3916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3881 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .X(net3917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3882 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[4] ),
    .X(net3918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3883 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[0] ),
    .X(net3919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3884 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ),
    .X(net3920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3885 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[2] ),
    .X(net3921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3886 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[2] ),
    .X(net3922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3887 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[2] ),
    .X(net3923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3888 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .X(net3924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3889 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[27] ),
    .X(net3925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3890 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[12] ),
    .X(net3926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3891 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .X(net3927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3892 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .X(net3928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3893 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ),
    .X(net3929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3894 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .X(net3930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3895 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .X(net3931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3896 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[7] ),
    .X(net3932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3897 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[10] ),
    .X(net3933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3898 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .X(net3934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3899 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[14] ),
    .X(net3935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3900 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .X(net3936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3901 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(net3937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3902 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[11] ),
    .X(net3938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3903 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .X(net3939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3904 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .X(net3940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3905 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[9] ),
    .X(net3941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3906 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[2] ),
    .X(net3942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3907 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .X(net3943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3908 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(net3944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3909 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[8] ),
    .X(net3945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3910 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[13] ),
    .X(net3946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3911 (.A(_04295_),
    .X(net3947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3912 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.o_[2] ),
    .X(net3948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3913 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .X(net3949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3914 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .X(net3950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3915 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[28] ),
    .X(net3951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3916 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[6] ),
    .X(net3952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3917 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(net3953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3918 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(net3954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3919 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[13] ),
    .X(net3955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3920 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(net3956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3921 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[0] ),
    .X(net3957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3922 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[3] ),
    .X(net3958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3923 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(net3959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3924 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .X(net3960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3925 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .X(net3961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3926 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(net3962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3927 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .X(net3963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3928 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[2] ),
    .X(net3964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3929 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(net3965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3930 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .X(net3966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3931 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(net3967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3932 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[31] ),
    .X(net3968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3933 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[3] ),
    .X(net3969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3934 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[35] ),
    .X(net3970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3935 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(net3971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3936 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(net3972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3937 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(net3973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3938 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[0] ),
    .X(net3974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3939 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(net3975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3940 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[6] ),
    .X(net3976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3941 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[36] ),
    .X(net3977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3942 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[39] ),
    .X(net3978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3943 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ),
    .X(net3979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3944 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(net3980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3945 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[3] ),
    .X(net3981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3946 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(net3982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3947 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[11] ),
    .X(net3983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3948 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[23] ),
    .X(net3984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3949 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .X(net3985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3950 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(net3986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3951 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[11] ),
    .X(net3987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3952 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(net3988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3953 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(net3989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3954 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[6] ),
    .X(net3990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3955 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(net3991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3956 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .X(net3992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3957 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[8] ),
    .X(net3993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3958 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[27] ),
    .X(net3994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3959 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[22] ),
    .X(net3995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3960 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[3] ),
    .X(net3996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3961 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[14] ),
    .X(net3997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3962 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[8] ),
    .X(net3998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3963 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[34] ),
    .X(net3999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3964 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .X(net4000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3965 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ),
    .X(net4001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3966 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(net4002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3967 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(net4003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3968 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[0] ),
    .X(net4004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3969 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(net4005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3970 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[23] ),
    .X(net4006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3971 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ),
    .X(net4007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3972 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ),
    .X(net4008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3973 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(net4009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3974 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ),
    .X(net4010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3975 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(net4011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3976 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[38] ),
    .X(net4012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3977 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(net4013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3978 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[6] ),
    .X(net4014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3979 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[11] ),
    .X(net4015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3980 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[30] ),
    .X(net4016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3981 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[1] ),
    .X(net4017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3982 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[1] ),
    .X(net4018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3983 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .X(net4019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3984 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(net4020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3985 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[3] ),
    .X(net4021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3986 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(net4022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3987 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[6] ),
    .X(net4023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3988 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .X(net4024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3989 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(net4025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3990 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[6] ),
    .X(net4026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3991 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[28] ),
    .X(net4027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3992 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[22] ),
    .X(net4028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3993 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .X(net4029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3994 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(net4030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3995 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .X(net4031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3996 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(net4032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3997 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[11] ),
    .X(net4033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3998 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(net4034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3999 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(net4035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4000 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(net4036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4001 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[8] ),
    .X(net4037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4002 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[27] ),
    .X(net4038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4003 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .X(net4039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4004 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ),
    .X(net4040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4005 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .X(net4041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4006 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[3] ),
    .X(net4042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4007 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ),
    .X(net4043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4008 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[6] ),
    .X(net4044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4009 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(net4045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4010 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .X(net4046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4011 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[20] ),
    .X(net4047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4012 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ),
    .X(net4048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4013 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(net4049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4014 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(net4050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4015 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[33] ),
    .X(net4051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4016 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .X(net4052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4017 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[11] ),
    .X(net4053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4018 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[15] ),
    .X(net4054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4019 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(net4055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4020 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(net4056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4021 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ),
    .X(net4057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4022 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.o[11] ),
    .X(net4058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4023 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .X(net4059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4024 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[9] ),
    .X(net4060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4025 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .X(net4061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4026 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ),
    .X(net4062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4027 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[17] ),
    .X(net4063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4028 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ),
    .X(net4064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4029 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[9] ),
    .X(net4065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4030 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[1] ),
    .X(net4066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4031 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(net4067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4032 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[7] ),
    .X(net4068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4033 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[37] ),
    .X(net4069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4034 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[25] ),
    .X(net4070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4035 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(net4071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4036 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[16] ),
    .X(net4072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4037 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[4] ),
    .X(net4073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4038 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(net4074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4039 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[8] ),
    .X(net4075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4040 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[4] ),
    .X(net4076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4041 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .X(net4077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4042 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[32] ),
    .X(net4078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4043 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[20] ),
    .X(net4079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4044 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[13] ),
    .X(net4080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4045 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .X(net4081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4046 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[3] ),
    .X(net4082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4047 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[7] ),
    .X(net4083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4048 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lb_in_sels[9] ),
    .X(net4084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4049 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[0] ),
    .X(net4085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4050 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ),
    .X(net4086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4051 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(net4087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4052 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(net4088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4053 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[3] ),
    .X(net4089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4054 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[12] ),
    .X(net4090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4055 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ),
    .X(net4091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4056 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[9] ),
    .X(net4092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4057 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(net4093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4058 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ),
    .X(net4094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4059 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[38] ),
    .X(net4095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4060 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ),
    .X(net4096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4061 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .X(net4097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4062 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[1] ),
    .X(net4098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4063 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[27] ),
    .X(net4099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4064 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[4] ),
    .X(net4100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4065 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .X(net4101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4066 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ),
    .X(net4102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4067 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[25] ),
    .X(net4103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4068 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ),
    .X(net4104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4069 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ),
    .X(net4105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4070 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[33] ),
    .X(net4106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4071 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ),
    .X(net4107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4072 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[26] ),
    .X(net4108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4073 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[8] ),
    .X(net4109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4074 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[4] ),
    .X(net4110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4075 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .X(net4111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4076 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ),
    .X(net4112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4077 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[36] ),
    .X(net4113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4078 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[25] ),
    .X(net4114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4079 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(net4115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4080 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .X(net4116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4081 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ),
    .X(net4117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4082 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ),
    .X(net4118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4083 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .X(net4119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4084 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[20] ),
    .X(net4120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4085 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .X(net4121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4086 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ),
    .X(net4122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4087 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[0] ),
    .X(net4123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4088 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[3] ),
    .X(net4124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4089 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .X(net4125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4090 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[0] ),
    .X(net4126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4091 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[9] ),
    .X(net4127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4092 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[15] ),
    .X(net4128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4093 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .X(net4129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4094 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[9] ),
    .X(net4130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4095 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ),
    .X(net4131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4096 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(net4132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4097 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[17] ),
    .X(net4133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4098 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ),
    .X(net4134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4099 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[15] ),
    .X(net4135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4100 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[7] ),
    .X(net4136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4101 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[12] ),
    .X(net4137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4102 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[30] ),
    .X(net4138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4103 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[28] ),
    .X(net4139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4104 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .X(net4140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4105 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(net4141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4106 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[2] ),
    .X(net4142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4107 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .X(net4143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4108 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ),
    .X(net4144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4109 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[10] ),
    .X(net4145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4110 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[3] ),
    .X(net4146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4111 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ),
    .X(net4147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4112 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ),
    .X(net4148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4113 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[4] ),
    .X(net4149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4114 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ),
    .X(net4150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4115 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.seg[1] ),
    .X(net4151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4116 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(net4152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4117 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[8] ),
    .X(net4153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4118 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .X(net4154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4119 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[0] ),
    .X(net4155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4120 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(net4156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4121 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ),
    .X(net4157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4122 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ),
    .X(net4158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4123 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[5] ),
    .X(net4159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4124 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(net4160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4125 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[8] ),
    .X(net4161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4126 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[1] ),
    .X(net4162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4127 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ),
    .X(net4163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4128 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[15] ),
    .X(net4164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4129 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ),
    .X(net4165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4130 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[26] ),
    .X(net4166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4131 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(net4167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4132 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ),
    .X(net4168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4133 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[3] ),
    .X(net4169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4134 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[3] ),
    .X(net4170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4135 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(net4171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4136 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[13] ),
    .X(net4172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4137 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[10] ),
    .X(net4173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4138 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ),
    .X(net4174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4139 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(net4175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4140 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[18] ),
    .X(net4176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4141 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[12] ),
    .X(net4177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4142 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ),
    .X(net4178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4143 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(net4179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4144 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[2] ),
    .X(net4180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4145 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ),
    .X(net4181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4146 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .X(net4182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4147 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.lut_in_sels[3] ),
    .X(net4183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4148 (.A(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ),
    .X(net4184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4149 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[15] ),
    .X(net4185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4150 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .X(net4186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4151 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[5] ),
    .X(net4187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4152 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[2] ),
    .X(net4188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4153 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.seg[3] ),
    .X(net4189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4154 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[10] ),
    .X(net4190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4155 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lb_in_sels[9] ),
    .X(net4191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4156 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ),
    .X(net4192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4157 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[16] ),
    .X(net4193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4158 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[13] ),
    .X(net4194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4159 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[0] ),
    .X(net4195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4160 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ),
    .X(net4196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4161 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[13] ),
    .X(net4197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4162 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[4] ),
    .X(net4198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4163 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(net4199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4164 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ),
    .X(net4200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4165 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[5] ),
    .X(net4201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4166 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[12] ),
    .X(net4202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4167 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ),
    .X(net4203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4168 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(net4204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4169 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ),
    .X(net4205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4170 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[8] ),
    .X(net4206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4171 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ),
    .X(net4207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4172 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[2] ),
    .X(net4208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4173 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[28] ),
    .X(net4209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4174 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.lut_in_sels[5] ),
    .X(net4210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4175 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[3] ),
    .X(net4211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4176 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ),
    .X(net4212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4177 (.A(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[9] ),
    .X(net4213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4178 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[34] ),
    .X(net4214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4179 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][16] ),
    .X(net4215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4180 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[0] ),
    .X(net4216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4181 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(net4217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4182 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.lb_in_sels[9] ),
    .X(net4218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4183 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.lb_in_sels[11] ),
    .X(net4219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4184 (.A(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(net4220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4185 (.A(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(net4221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4186 (.A(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.seg[0] ),
    .X(net4222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4187 (.A(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.seg[1] ),
    .X(net4223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4188 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[23] ),
    .X(net4224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4189 (.A(_04045_),
    .X(net4225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4190 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.o_[4] ),
    .X(net4226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4191 (.A(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(net4227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4192 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.seg[0] ),
    .X(net4228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4193 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.luts.seg[0] ),
    .X(net4229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4194 (.A(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.luts.seg[0] ),
    .X(net4230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4195 (.A(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[13] ),
    .X(net4231));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__A (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__A (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__A (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__A (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06303__A (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05330__A (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05171__A (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05017__A (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04887__A (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04815__A (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08784__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06822__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06387__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05304__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04816__A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__A0 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__A0 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__A0 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10020__A0 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__A0 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05494__A1 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05485__A1 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05476__A1 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05280__A1 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04827__A1 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08198__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05278__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04930__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04888__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04877__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04870__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04863__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04825__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__B1 (.DIODE(_00181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06931__A (.DIODE(_00181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06669__A (.DIODE(_00181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05532__B1 (.DIODE(_00181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05511__B1 (.DIODE(_00181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05502__B1 (.DIODE(_00181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05466__B1 (.DIODE(_00181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05062__A (.DIODE(_00181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04880__A (.DIODE(_00181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04826__B1 (.DIODE(_00181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06393__A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05314__A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04918__A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04830__A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__A0 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__A0 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A0 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A0 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__A0 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05496__A1 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05487__A1 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05478__A1 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05282__A1 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04831__A1 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06315__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05341__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05317__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05182__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05028__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04908__B (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04834__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06759__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05527__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04973__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04835__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10119__A0 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__A0 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__A0 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__A0 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__A0 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05498__A1 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05489__A1 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05480__A1 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05284__A1 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04836__A1 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06282__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04976__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04839__A (.DIODE(_00191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10121__A0 (.DIODE(_00192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10111__A0 (.DIODE(_00192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A0 (.DIODE(_00192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__A0 (.DIODE(_00192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__A0 (.DIODE(_00192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__A0 (.DIODE(_00192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__A0 (.DIODE(_00192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__A0 (.DIODE(_00192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__A0 (.DIODE(_00192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04840__A1 (.DIODE(_00192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A (.DIODE(_00195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__A (.DIODE(_00195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09578__A (.DIODE(_00195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A (.DIODE(_00195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08687__A (.DIODE(_00195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A (.DIODE(_00195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A (.DIODE(_00195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04966__B1 (.DIODE(_00195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04874__A (.DIODE(_00195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04844__A (.DIODE(_00195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10651__A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06855__A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05379__A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05067__A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04948__A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04845__A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04947__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04940__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04938__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04936__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04904__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04895__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04893__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04873__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04866__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04859__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__C1 (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__C1 (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__C1 (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__C1 (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__C1 (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__C1 (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__C1 (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__C1 (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__C1 (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04858__A (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06309__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05225__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05071__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04957__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04947__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04936__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04917__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04859__B1 (.DIODE(_00210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05337__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05178__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05024__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04861__A (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__A (.DIODE(_00215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A (.DIODE(_00215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A (.DIODE(_00215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__A (.DIODE(_00215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05228__A (.DIODE(_00215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04865__A (.DIODE(_00215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05088__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05074__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04959__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04950__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04938__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04921__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04904__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04893__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04866__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04990__A2 (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04922__A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04906__A1 (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04868__A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__C1 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__C1 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__C1 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__C1 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__C1 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__A (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__A (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05104__A (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04924__A (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04872__A (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06365__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06317__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04961__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04952__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04940__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04895__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04873__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__A1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__A1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04963__A1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04954__A1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04925__A1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04921__A1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04917__A1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04913__A1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04897__A1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04879__A1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__A (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__A (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__A (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05408__A (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04943__A (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04878__A (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__B1 (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05148__A (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04963__B1_N (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04954__B1_N (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04926__A (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04913__B1_N (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04897__B1_N (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04879__B1_N (.DIODE(_00227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__B1 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__B1 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__C1 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10074__C1 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__C1 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__C1 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__C1 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__C1 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05023__A (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04881__A (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__A (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05022__A1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04994__A1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04991__A1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04988__A1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04983__A1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04944__A1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04911__A1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04902__A1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04891__A1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04896__S (.DIODE(_00233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04894__S (.DIODE(_00233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04892__S (.DIODE(_00233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04886__S (.DIODE(_00233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__A1 (.DIODE(_00235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__A1 (.DIODE(_00235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__A1 (.DIODE(_00235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__A1 (.DIODE(_00235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__A (.DIODE(_00235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A (.DIODE(_00235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__A (.DIODE(_00235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05520__A (.DIODE(_00235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04964__A (.DIODE(_00235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04889__A (.DIODE(_00235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10562__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06346__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04986__A (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04889__B (.DIODE(_00236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10125__B1 (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__B1 (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10039__B1 (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05398__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05176__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04890__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05139__B1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05112__B1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05098__B1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05085__B1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05055__B1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05041__B1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05022__B1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04983__B1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04902__B1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04891__B1 (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__B1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10076__B1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__B1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__B1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__B1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__B1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__B1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09195__B1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04908__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__B1 (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10047__B1 (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__B1 (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__B1 (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__B1 (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__B1 (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__B1 (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06838__A (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05217__A (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04910__A (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05203__B1 (.DIODE(_00252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05185__B1 (.DIODE(_00252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05145__B1 (.DIODE(_00252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05118__B1 (.DIODE(_00252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05091__B1 (.DIODE(_00252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05061__B1 (.DIODE(_00252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05047__B1 (.DIODE(_00252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05031__B1 (.DIODE(_00252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04991__B1 (.DIODE(_00252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04911__B1 (.DIODE(_00252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__B1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__B1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__B1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__B1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__B1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__B1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__B1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__B1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05077__B1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04925__B1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06869__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06348__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05435__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05393__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05277__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05235__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05121__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05080__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04933__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08834__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05345__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05186__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05032__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04928__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__B1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__B1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__B1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06846__B1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06325__B1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05311__B1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05157__B1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05003__B1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04931__A (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__A (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__A (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__A (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05434__C1 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05392__C1 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05276__C1 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05234__C1 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05120__C1 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05079__C1 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04932__C1 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__A (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__A (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__A (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05108__B1 (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05094__B1 (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05066__B1 (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05050__B1 (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05035__B1 (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04994__B1 (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04944__B1 (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06365__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06317__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06309__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04961__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04959__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04957__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04952__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04950__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__A1 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__A1 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__A1 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__A1 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A1 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A1 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05158__A0 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05126__A0 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05004__A0 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04967__A0 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__A1 (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__A1 (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__A1 (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__A1 (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__A (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__A (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__A (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05524__A (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04986__B (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04970__A (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05160__A0 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05128__A0 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05006__A0 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04971__A0 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A1 (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__A1 (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A1 (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__A1 (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__A1 (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__A1 (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05162__A0 (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05130__A0 (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05008__A0 (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04974__A0 (.DIODE(_00295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05539__A0 (.DIODE(_00297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05518__A0 (.DIODE(_00297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05509__A0 (.DIODE(_00297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05473__A0 (.DIODE(_00297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05444__A0 (.DIODE(_00297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05321__A0 (.DIODE(_00297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05164__A0 (.DIODE(_00297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05132__A0 (.DIODE(_00297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05010__A0 (.DIODE(_00297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04977__A0 (.DIODE(_00297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__B1 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__B1 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08828__A (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06362__A (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05257__A (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04987__A (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05214__B1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05199__B1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05181__B1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05142__B1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05115__B1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05101__B1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05058__B1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05044__B1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05027__B1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04988__B1 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__A (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05463__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05305__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04996__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05038__C_N (.DIODE(_00312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04997__A (.DIODE(_00312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05138__A2 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05111__A1 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05097__A1 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05084__A1 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05069__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05054__A1 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05040__A0 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05021__A3 (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__B1 (.DIODE(_00332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__B1 (.DIODE(_00332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05021__B2 (.DIODE(_00332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05061__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05058__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05055__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05050__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05047__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05044__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05041__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05035__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05031__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05027__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05141__A2 (.DIODE(_00335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05114__A1 (.DIODE(_00335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05100__A1 (.DIODE(_00335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05087__A (.DIODE(_00335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05072__A (.DIODE(_00335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05057__A1 (.DIODE(_00335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05043__A0 (.DIODE(_00335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05026__A3 (.DIODE(_00335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__S1 (.DIODE(_00336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05026__B2 (.DIODE(_00336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05144__A2 (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05117__A1 (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05102__A (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05090__A1 (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05075__A (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05060__A1 (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05046__A0 (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05030__A3 (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__A (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__A (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06830__A (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05446__A (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05375__A (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05336__A (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05254__A (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05200__A (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05134__A (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05063__A (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__S1 (.DIODE(_00365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05065__A0 (.DIODE(_00365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05261__A1 (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05243__A1 (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05232__A1 (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05229__A1 (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05225__A1 (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05105__A1 (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05088__A1 (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05077__A1 (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05074__A1 (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05071__A1 (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__B1 (.DIODE(_00394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__B1 (.DIODE(_00394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__B1 (.DIODE(_00394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06866__B1 (.DIODE(_00394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06344__B1 (.DIODE(_00394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05419__B1 (.DIODE(_00394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05390__B1 (.DIODE(_00394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05261__B1 (.DIODE(_00394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05232__B1 (.DIODE(_00394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05105__B1 (.DIODE(_00394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__B1 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09569__B1 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__B1 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__B1 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B1 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08301__A (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06377__A (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05124__A (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07095__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06289__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06275__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05437__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05125__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05132__S (.DIODE(_00409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05130__S (.DIODE(_00409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05128__S (.DIODE(_00409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05126__S (.DIODE(_00409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05199__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05196__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05189__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05185__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05181__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05177__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05149__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05145__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05142__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05139__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05378__B1 (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05363__B1 (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05348__B1 (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05303__B1 (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05264__B1 (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05249__B1 (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05221__B1 (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05206__B1 (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05189__B1 (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05149__B1 (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05164__S (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05162__S (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05160__S (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05158__S (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05293__A2 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05267__A1 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05252__A1 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05239__A1 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05223__A (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05210__A1 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05195__A0 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05175__A3 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09728__B1 (.DIODE(_00446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05175__B2 (.DIODE(_00446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05368__B1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05354__B1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05335__B1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05294__B1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05268__B1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05253__B1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05240__B1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05211__B1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05196__B1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05177__B1 (.DIODE(_00448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05296__A2 (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05270__A1 (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05256__A1 (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05242__A (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05226__A (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05213__A1 (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05198__A0 (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05180__A3 (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05302__A2 (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05276__A1 (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05263__A1 (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05248__A1 (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05234__A1 (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05220__A1 (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05205__A0 (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05188__A3 (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05253__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05249__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05246__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05240__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05221__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05218__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05214__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05211__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05206__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05203__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05220__S (.DIODE(_00473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05216__S (.DIODE(_00473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05213__S (.DIODE(_00473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05210__S (.DIODE(_00473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05457__B1 (.DIODE(_00479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05432__B1 (.DIODE(_00479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05405__B1 (.DIODE(_00479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05374__B1 (.DIODE(_00479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05360__B1 (.DIODE(_00479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05344__B1 (.DIODE(_00479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05300__B1 (.DIODE(_00479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05274__B1 (.DIODE(_00479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05246__B1 (.DIODE(_00479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05218__B1 (.DIODE(_00479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05234__A2 (.DIODE(_00482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05233__B (.DIODE(_00482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05231__B (.DIODE(_00482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05230__B (.DIODE(_00482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05227__B (.DIODE(_00482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05226__B (.DIODE(_00482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05224__B (.DIODE(_00482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05223__B (.DIODE(_00482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__B1 (.DIODE(_00487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07010__B1 (.DIODE(_00487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06923__B1 (.DIODE(_00487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__B1 (.DIODE(_00487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06576__B1 (.DIODE(_00487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06341__B1 (.DIODE(_00487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05402__B1 (.DIODE(_00487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05387__B1 (.DIODE(_00487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05243__B1 (.DIODE(_00487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05229__B1 (.DIODE(_00487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05248__S (.DIODE(_00494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05245__S (.DIODE(_00494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05242__B (.DIODE(_00494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05241__B (.DIODE(_00494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05239__S (.DIODE(_00494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05263__S (.DIODE(_00503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05260__B (.DIODE(_00503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05259__B (.DIODE(_00503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05256__S (.DIODE(_00503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05252__S (.DIODE(_00503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05335__A1 (.DIODE(_00505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05303__A1 (.DIODE(_00505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05300__A1 (.DIODE(_00505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05297__A1 (.DIODE(_00505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05294__A1 (.DIODE(_00505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05274__A1 (.DIODE(_00505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05271__A1 (.DIODE(_00505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05268__A1 (.DIODE(_00505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05264__A1 (.DIODE(_00505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05258__A1 (.DIODE(_00505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06314__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05454__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05429__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05416__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05371__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05357__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05340__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05297__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05271__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05258__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05276__A2 (.DIODE(_00514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05275__B (.DIODE(_00514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05273__S (.DIODE(_00514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05270__S (.DIODE(_00514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05267__S (.DIODE(_00514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06368__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06349__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05521__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05493__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05484__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05475__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05279__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__A1 (.DIODE(_00527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A1 (.DIODE(_00527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09830__A1 (.DIODE(_00527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__A1 (.DIODE(_00527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09556__A1 (.DIODE(_00527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__A1 (.DIODE(_00527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__A1 (.DIODE(_00527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__A1 (.DIODE(_00527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__A (.DIODE(_00527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05287__A (.DIODE(_00527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__A1 (.DIODE(_00528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__A1 (.DIODE(_00528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__A1 (.DIODE(_00528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06375__A1 (.DIODE(_00528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06356__A1 (.DIODE(_00528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05530__A1 (.DIODE(_00528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05500__A1 (.DIODE(_00528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05491__A1 (.DIODE(_00528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05482__A1 (.DIODE(_00528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05288__A1 (.DIODE(_00528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06379__A0 (.DIODE(_00540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06326__A0 (.DIODE(_00540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06290__A0 (.DIODE(_00540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06276__A0 (.DIODE(_00540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05533__A0 (.DIODE(_00540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05512__A0 (.DIODE(_00540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05503__A0 (.DIODE(_00540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05467__A0 (.DIODE(_00540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05438__A0 (.DIODE(_00540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05312__A0 (.DIODE(_00540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06381__A0 (.DIODE(_00549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06328__A0 (.DIODE(_00549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06292__A0 (.DIODE(_00549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06278__A0 (.DIODE(_00549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05535__A0 (.DIODE(_00549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05514__A0 (.DIODE(_00549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05505__A0 (.DIODE(_00549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05469__A0 (.DIODE(_00549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05440__A0 (.DIODE(_00549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05315__A0 (.DIODE(_00549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A (.DIODE(_00551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__A (.DIODE(_00551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08456__A (.DIODE(_00551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__A (.DIODE(_00551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__A (.DIODE(_00551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__A (.DIODE(_00551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__A (.DIODE(_00551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06836__A (.DIODE(_00551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06476__A (.DIODE(_00551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05318__A (.DIODE(_00551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06383__A0 (.DIODE(_00552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06330__A0 (.DIODE(_00552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06294__A0 (.DIODE(_00552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06280__A0 (.DIODE(_00552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05537__A0 (.DIODE(_00552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05516__A0 (.DIODE(_00552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05507__A0 (.DIODE(_00552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05471__A0 (.DIODE(_00552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05442__A0 (.DIODE(_00552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05319__A0 (.DIODE(_00552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05453__A2 (.DIODE(_00568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05428__A1 (.DIODE(_00568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05415__A1 (.DIODE(_00568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05401__A (.DIODE(_00568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05385__A (.DIODE(_00568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05370__A1 (.DIODE(_00568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05356__A0 (.DIODE(_00568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05339__A3 (.DIODE(_00568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__S1 (.DIODE(_00569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05339__B2 (.DIODE(_00569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05459__A2 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05434__A1 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05421__A1 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05407__A1 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05392__A1 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05377__A1 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05362__A0 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05347__A3 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05432__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05429__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05426__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05422__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05416__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05413__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05409__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05405__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05399__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05378__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06576__A1 (.DIODE(_00599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06494__A1 (.DIODE(_00599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06344__A1 (.DIODE(_00599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06341__A1 (.DIODE(_00599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06338__A1 (.DIODE(_00599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05419__A1 (.DIODE(_00599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05402__A1 (.DIODE(_00599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05390__A1 (.DIODE(_00599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05387__A1 (.DIODE(_00599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05384__A1 (.DIODE(_00599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__B1 (.DIODE(_00603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__B1 (.DIODE(_00603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__B1 (.DIODE(_00603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__B1 (.DIODE(_00603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__B1 (.DIODE(_00603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__B1 (.DIODE(_00603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__B1 (.DIODE(_00603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06494__B1 (.DIODE(_00603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06338__B1 (.DIODE(_00603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05384__B1 (.DIODE(_00603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__B1 (.DIODE(_00614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__B1 (.DIODE(_00614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__B1 (.DIODE(_00614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06881__B1 (.DIODE(_00614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__B1 (.DIODE(_00614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06360__B1 (.DIODE(_00614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05451__B1 (.DIODE(_00614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05426__B1 (.DIODE(_00614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05413__B1 (.DIODE(_00614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05399__B1 (.DIODE(_00614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__B1 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__B1 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06929__B1 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06887__B1 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06843__B1 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06367__B1 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06322__B1 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05460__B1 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05422__B1 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05409__B1 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__A1 (.DIODE(_00646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06367__A1 (.DIODE(_00646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06363__A1 (.DIODE(_00646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06360__A1 (.DIODE(_00646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06322__A1 (.DIODE(_00646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06314__A1 (.DIODE(_00646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05460__A1 (.DIODE(_00646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05457__A1 (.DIODE(_00646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05454__A1 (.DIODE(_00646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05451__A1 (.DIODE(_00646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05473__S (.DIODE(_00662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05471__S (.DIODE(_00662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05469__S (.DIODE(_00662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05467__S (.DIODE(_00662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05482__S (.DIODE(_00667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05480__S (.DIODE(_00667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05478__S (.DIODE(_00667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05476__S (.DIODE(_00667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05491__S (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05489__S (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05487__S (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05485__S (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05500__S (.DIODE(_00677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05498__S (.DIODE(_00677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05496__S (.DIODE(_00677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05494__S (.DIODE(_00677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05509__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05507__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05505__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05503__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A1 (.DIODE(_00692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__A1 (.DIODE(_00692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A1 (.DIODE(_00692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__A1 (.DIODE(_00692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__A1 (.DIODE(_00692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__A1 (.DIODE(_00692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__A1 (.DIODE(_00692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06369__A1 (.DIODE(_00692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06350__A1 (.DIODE(_00692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05522__A1 (.DIODE(_00692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05530__S (.DIODE(_00693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05528__S (.DIODE(_00693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05525__S (.DIODE(_00693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05522__S (.DIODE(_00693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__A1 (.DIODE(_00695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__A1 (.DIODE(_00695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__A1 (.DIODE(_00695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__A1 (.DIODE(_00695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__A1 (.DIODE(_00695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__A1 (.DIODE(_00695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__A1 (.DIODE(_00695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06371__A1 (.DIODE(_00695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06352__A1 (.DIODE(_00695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05525__A1 (.DIODE(_00695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07024__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06373__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06354__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05528__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06472__A (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06158__C1 (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05986__C1 (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05808__C1 (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05619__C1 (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05620__B2 (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__A0 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__A0 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__A0 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08770__A0 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__A0 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05627__A0 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05621__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__A3 (.DIODE(_00788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A0 (.DIODE(_00788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__A2 (.DIODE(_00788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08760__A2 (.DIODE(_00788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__A2 (.DIODE(_00788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A2 (.DIODE(_00788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A0 (.DIODE(_00788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05990__A2 (.DIODE(_00788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05905__A2 (.DIODE(_00788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05627__A2 (.DIODE(_00788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__B (.DIODE(_00792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A2 (.DIODE(_00792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__A2 (.DIODE(_00792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__A2 (.DIODE(_00792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__A2 (.DIODE(_00792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__A2 (.DIODE(_00792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A2 (.DIODE(_00792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A1 (.DIODE(_00792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06079__A2 (.DIODE(_00792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05631__A2 (.DIODE(_00792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__B (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08762__A3 (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__A3 (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A3 (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A3 (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A3 (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06079__A3 (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05992__A3 (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05907__A3 (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05631__A3 (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__B2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05711__B2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05707__B1 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05701__A (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05678__A (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05709__S (.DIODE(_00824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05708__S (.DIODE(_00824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05706__S (.DIODE(_00824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05702__S (.DIODE(_00824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05699__S (.DIODE(_00824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05698__S (.DIODE(_00824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05664__S (.DIODE(_00824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05663__S (.DIODE(_00824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05710__S (.DIODE(_00838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05707__A1 (.DIODE(_00838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05703__A (.DIODE(_00838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05700__S (.DIODE(_00838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05677__S (.DIODE(_00838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05712__A2 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05711__C1 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05717__A2 (.DIODE(_00874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__A (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__A0 (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__A0 (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05719__A (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05718__A (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__A0 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A0 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A0 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__A0 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A0 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__A0 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__A (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__A0 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06251__A0 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05723__A0 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A1 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__A2 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__A0 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__A2 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A0 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06265__A1 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__A2 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06253__A0 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05815__A2 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__A0 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__A3 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__A1 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__A3 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A1 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06262__A1 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__A3 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06253__A1 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06162__A1 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05815__A3 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__A1 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__B (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A2 (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06265__A2 (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06262__A2 (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06257__A2 (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06253__A2 (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__A2 (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06162__A2 (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05818__A2 (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__A2 (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__B (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A3 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06265__A3 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06262__A3 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06257__A3 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06253__A3 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__A3 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06162__A3 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05818__A3 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__A3 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__A1 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__A1 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05812__A1 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05805__S (.DIODE(_00938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05802__A1 (.DIODE(_00938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05800__B1 (.DIODE(_00938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05782__S (.DIODE(_00938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05779__S (.DIODE(_00938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__A2 (.DIODE(_00968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__A2 (.DIODE(_00968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05812__A2 (.DIODE(_00968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__C1 (.DIODE(_00971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__C1 (.DIODE(_00971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05812__B1 (.DIODE(_00971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A1 (.DIODE(_00972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__A (.DIODE(_00972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__A1 (.DIODE(_00972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A1 (.DIODE(_00972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__A1 (.DIODE(_00972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__A (.DIODE(_00972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__A1 (.DIODE(_00972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05813__A (.DIODE(_00972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A3 (.DIODE(_00973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A3 (.DIODE(_00973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A1 (.DIODE(_00973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__A1 (.DIODE(_00973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06267__A3 (.DIODE(_00973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06261__A3 (.DIODE(_00973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__A1 (.DIODE(_00973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06247__A1 (.DIODE(_00973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06161__A1 (.DIODE(_00973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05815__A1 (.DIODE(_00973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A0 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A0 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A0 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A0 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06267__A0 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06261__A0 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06257__A0 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06247__A2 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06161__A2 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05818__A0 (.DIODE(_00975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A1 (.DIODE(_00976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A3 (.DIODE(_00976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A3 (.DIODE(_00976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A1 (.DIODE(_00976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06267__A1 (.DIODE(_00976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06261__A1 (.DIODE(_00976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06257__A1 (.DIODE(_00976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06247__A3 (.DIODE(_00976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06161__A3 (.DIODE(_00976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05818__A1 (.DIODE(_00976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05895__A2 (.DIODE(_01007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05894__B (.DIODE(_01007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05891__S (.DIODE(_01007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05889__S (.DIODE(_01007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05888__S (.DIODE(_01007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05867__S (.DIODE(_01007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05866__S (.DIODE(_01007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05851__S (.DIODE(_01007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05850__S (.DIODE(_01007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05895__B1 (.DIODE(_01020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05892__A1 (.DIODE(_01020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05890__S (.DIODE(_01020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05868__S (.DIODE(_01020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05863__S (.DIODE(_01020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05898__B2 (.DIODE(_01055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__A3 (.DIODE(_01056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__A3 (.DIODE(_01056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A (.DIODE(_01056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__A1 (.DIODE(_01056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__A0 (.DIODE(_01056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A0 (.DIODE(_01056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05905__A0 (.DIODE(_01056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05899__A (.DIODE(_01056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08946__A2 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__A0 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A3 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__A2 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__A2 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A1 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A3 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06077__A2 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05990__A1 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05905__A1 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A1 (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A1 (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05904__A (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08946__A3 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__A2 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__A3 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__A3 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08760__A3 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__A3 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A3 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06077__A3 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05990__A3 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05905__A3 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05987__B2 (.DIODE(_01142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__A1 (.DIODE(_01143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__A1 (.DIODE(_01143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__A (.DIODE(_01143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A2 (.DIODE(_01143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08760__A0 (.DIODE(_01143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A2 (.DIODE(_01143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05990__A0 (.DIODE(_01143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05988__A (.DIODE(_01143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06069__S (.DIODE(_01176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06065__S (.DIODE(_01176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06063__S (.DIODE(_01176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06062__S (.DIODE(_01176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06059__S (.DIODE(_01176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06058__S (.DIODE(_01176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06024__S (.DIODE(_01176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06023__S (.DIODE(_01176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06070__A1 (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06066__A (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06064__S (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06060__S (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06037__S (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06073__B2 (.DIODE(_01226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__A2 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__A2 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__A (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08946__A0 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__A0 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__A0 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06077__A0 (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06074__A (.DIODE(_01227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06159__B2 (.DIODE(_01310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__A (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A2 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__A2 (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__A (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08965__A (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06160__A (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06241__S (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06240__A2 (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06239__A_N (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06237__S (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06234__S (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06210__S (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06209__S (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06195__S (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06194__S (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06768__B2 (.DIODE(_01356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06242__B2 (.DIODE(_01356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06238__S (.DIODE(_01356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06211__S (.DIODE(_01356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06207__S (.DIODE(_01356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06245__B2 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09336__A (.DIODE(_01395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A3 (.DIODE(_01395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__A3 (.DIODE(_01395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09026__A (.DIODE(_01395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__A (.DIODE(_01395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06246__A (.DIODE(_01395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__C (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09420__C (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__B (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__B (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__B (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__C (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__C (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__C (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06298__B (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06272__B (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__A0 (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__A0 (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06853__A0 (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__A0 (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06806__A0 (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06479__A0 (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06385__A0 (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06332__A0 (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06296__A0 (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06283__A0 (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06493__A (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06359__A1 (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06336__A (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06304__B (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10040__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07655__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06832__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06312__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06574__A (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06361__A1 (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06339__A (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06313__A1 (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09149__A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06841__A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06320__A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__C1 (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__C1 (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__C1 (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__C1 (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__C1 (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__C1 (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__C1 (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06868__C1 (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__C1 (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06347__C1 (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06356__S (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06354__S (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06352__S (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06350__S (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__B1 (.DIODE(_01481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__B1 (.DIODE(_01481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__B1 (.DIODE(_01481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__B1 (.DIODE(_01481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__B1 (.DIODE(_01481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__B1 (.DIODE(_01481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__B1 (.DIODE(_01481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__B1 (.DIODE(_01481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06834__B1 (.DIODE(_01481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06363__B1 (.DIODE(_01481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06375__S (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06373__S (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06371__S (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06369__S (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__B1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__B1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09746__B1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__B1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09439__B1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__B1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__B1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__B1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__B1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06378__B1 (.DIODE(_01489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__A0 (.DIODE(_01495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__A0 (.DIODE(_01495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A0 (.DIODE(_01495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__A0 (.DIODE(_01495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06909__A0 (.DIODE(_01495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__A0 (.DIODE(_01495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__A0 (.DIODE(_01495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__A0 (.DIODE(_01495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__A0 (.DIODE(_01495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06391__A0 (.DIODE(_01495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__B1 (.DIODE(_01497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__B1 (.DIODE(_01497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__B1 (.DIODE(_01497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__B1 (.DIODE(_01497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__B1 (.DIODE(_01497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B1 (.DIODE(_01497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__B1 (.DIODE(_01497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__B1 (.DIODE(_01497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06908__B1 (.DIODE(_01497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06390__B1 (.DIODE(_01497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A0 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A0 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__A0 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__A0 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06911__A0 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__A0 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__A0 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__A0 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06802__A0 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06394__A0 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__A (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__A (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__C1 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__C1 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__C1 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06769__A (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__C1 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06661__C1 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06473__C1 (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06474__B2 (.DIODE(_01579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A0 (.DIODE(_01580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A0 (.DIODE(_01580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__A (.DIODE(_01580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09004__A (.DIODE(_01580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__A (.DIODE(_01580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06475__A (.DIODE(_01580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A0 (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__A0 (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A0 (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__A0 (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__A0 (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__A0 (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__A0 (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__A0 (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__A0 (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06477__A0 (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A0 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A0 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A0 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A0 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A0 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__A0 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__A2 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__A0 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06675__A0 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__A2 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A3 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__A3 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A3 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A3 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__A3 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__A3 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__A3 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06763__A1 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06674__A1 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__A3 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A2 (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A0 (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A2 (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A0 (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A1 (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__A2 (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__A0 (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__A1 (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06578__A2 (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__A0 (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A3 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A1 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A3 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A1 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__A1 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__A3 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__A1 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06675__A1 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06578__A3 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__A1 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__B (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A2 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A2 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__A2 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__A2 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__A2 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__A2 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06675__A2 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__A2 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__A2 (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__B (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A3 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A3 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__A3 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__A3 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__A3 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__A3 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06675__A3 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__A3 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__A3 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06572__B2 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A1 (.DIODE(_01673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A1 (.DIODE(_01673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__A (.DIODE(_01673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__A (.DIODE(_01673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__A (.DIODE(_01673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06573__A (.DIODE(_01673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__A1 (.DIODE(_01676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A1 (.DIODE(_01676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A3 (.DIODE(_01676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A3 (.DIODE(_01676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A1 (.DIODE(_01676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__A1 (.DIODE(_01676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__A1 (.DIODE(_01676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06763__A3 (.DIODE(_01676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06674__A3 (.DIODE(_01676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06578__A1 (.DIODE(_01676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__A2 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__A0 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A0 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A0 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A0 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__A2 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__A0 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06763__A0 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06674__A0 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__A0 (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06662__B2 (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09877__A (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09006__A (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__A (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06663__A (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__A1 (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__A1 (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A1 (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__A1 (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A1 (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__A1 (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__A1 (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__A1 (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__A1 (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__A1 (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__A2 (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__A2 (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__A2 (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06670__B (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09820__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08872__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08486__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06670__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__B1 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__B1 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__B1 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__C1 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__C1 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__C1 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__C1 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__C1 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__C1 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__C1 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10069__B1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__B1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09796__B1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__B1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__C1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__C1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__C1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__C1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__C1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__C1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__S (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06750__S (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06748__S (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06747__S (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06729__S (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06728__S (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06715__S (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__S (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06757__B2 (.DIODE(_01848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A3 (.DIODE(_01849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A3 (.DIODE(_01849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__A (.DIODE(_01849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09007__A (.DIODE(_01849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08956__A (.DIODE(_01849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06758__A (.DIODE(_01849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10132__B1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__B1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__B1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__B1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09191__B1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08920__B1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__B1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__B1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08690__B1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__C1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09296__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07088__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06770__B1 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__B (.DIODE(_01860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__A (.DIODE(_01862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__A (.DIODE(_01862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__S (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__S (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__S (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__S (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__S (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__S (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__S (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__S (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06939__S (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__S (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__C (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__C (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__C (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__C (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__C (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__C (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__B (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__C (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__C (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06795__C (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06806__S (.DIODE(_01883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__S (.DIODE(_01883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06802__S (.DIODE(_01883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__S (.DIODE(_01883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__B1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__B1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__B1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__B1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__B1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__B1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__B1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__B1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__B1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06839__B1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06853__S (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__S (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__S (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__S (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07010__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06923__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06866__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__A1 (.DIODE(_01923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__S (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__S (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__S (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__S (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__S (.DIODE(_01944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__S (.DIODE(_01944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__S (.DIODE(_01944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__S (.DIODE(_01944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__A2 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__A2 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__A2 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__B (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07084__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__C1 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__C1 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__C1 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__C1 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__C1 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__C1 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__C1 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__C1 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__C1 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__C1 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__S (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__S (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__S (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__S (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__A0 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A0 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A0 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__A0 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__A0 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07069__A0 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__A0 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__A0 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__A0 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__A0 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__S (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__S (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__S (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__S (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A (.DIODE(_02003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__A (.DIODE(_02003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A (.DIODE(_02003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A (.DIODE(_02003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__A (.DIODE(_02003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A (.DIODE(_02003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__A (.DIODE(_02003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__A (.DIODE(_02003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__A (.DIODE(_02003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__A (.DIODE(_02003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__S (.DIODE(_02019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__S (.DIODE(_02019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__S (.DIODE(_02019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__S (.DIODE(_02019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08358__A (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08197__A (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__A (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__A (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__A (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__A (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__A (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__A (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07017__A (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__B1 (.DIODE(_02034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08021__B1 (.DIODE(_02034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__B1 (.DIODE(_02034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07847__B1 (.DIODE(_02034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__B1 (.DIODE(_02034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__B1 (.DIODE(_02034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__B1 (.DIODE(_02034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__B1 (.DIODE(_02034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__B1 (.DIODE(_02034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__B1 (.DIODE(_02034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__S (.DIODE(_02035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07024__S (.DIODE(_02035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__S (.DIODE(_02035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__S (.DIODE(_02035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__A1 (.DIODE(_02044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__A1 (.DIODE(_02044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A1 (.DIODE(_02044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__A1 (.DIODE(_02044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__A1 (.DIODE(_02044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__A1 (.DIODE(_02044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__A1 (.DIODE(_02044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A1 (.DIODE(_02044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A1 (.DIODE(_02044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A1 (.DIODE(_02044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__S (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__S (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__S (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__S (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07854__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__A0 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A0 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__A0 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__A0 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__A0 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07556__A0 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__A0 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A0 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__A0 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__A0 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__A0 (.DIODE(_02062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A0 (.DIODE(_02062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A0 (.DIODE(_02062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__A0 (.DIODE(_02062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A0 (.DIODE(_02062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A0 (.DIODE(_02062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__A0 (.DIODE(_02062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__A0 (.DIODE(_02062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__A0 (.DIODE(_02062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07064__A0 (.DIODE(_02062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__A0 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__A0 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__A0 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__A0 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A0 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__A0 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A0 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__A0 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A0 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07067__A0 (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__A2 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__A2 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__A2 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07084__B (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__S (.DIODE(_02083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__S (.DIODE(_02083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__S (.DIODE(_02083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__S (.DIODE(_02083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__B1 (.DIODE(_02092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__B1 (.DIODE(_02092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__B1 (.DIODE(_02092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__B1 (.DIODE(_02092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__B1 (.DIODE(_02092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B1 (.DIODE(_02092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__B1 (.DIODE(_02092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07634__B1 (.DIODE(_02092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__B1 (.DIODE(_02092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07109__B1 (.DIODE(_02092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__S (.DIODE(_02093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__S (.DIODE(_02093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__S (.DIODE(_02093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__S (.DIODE(_02093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__S (.DIODE(_02121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__S (.DIODE(_02121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__S (.DIODE(_02121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__S (.DIODE(_02121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__A1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__A1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__A1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__A1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__A1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__A1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__S (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__S (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__S (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__S (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__B1 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08159__B1 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__B1 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07975__B1 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__B1 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__B1 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__B1 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07654__B1 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__B1 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__B1 (.DIODE(_02145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__A1 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A1 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__A1 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07654__A1 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__A1 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__A1 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__A1 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A1 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__A1 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__A1 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__S (.DIODE(_02191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__S (.DIODE(_02191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__S (.DIODE(_02191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__S (.DIODE(_02191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A0 (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__A0 (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A0 (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A0 (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__A0 (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__A0 (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__A0 (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__A (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08970__A (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__A (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A0 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A0 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__A0 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__A0 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A0 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__A0 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A2 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A0 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A0 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A2 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A3 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A3 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A1 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A3 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A3 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__A3 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A3 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A3 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A3 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A3 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A2 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__A0 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A2 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A0 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A1 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A2 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__A0 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A1 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A2 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A0 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A3 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__A1 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A3 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A1 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__A1 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A3 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__A1 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A1 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A3 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A1 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__B (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A2 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A2 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__A2 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__A2 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__A2 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A2 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A2 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A2 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A2 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__B (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A3 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A3 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__A3 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__A3 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__A3 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A3 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A3 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A3 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A3 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__B2 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09018__A (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__A3 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A3 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A3 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__A1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__A0 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A0 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A0 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A0 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A0 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__A2 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__A0 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A2 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A2 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A0 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__B2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A2 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__A2 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A2 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A2 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__A2 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__A2 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__A2 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__S (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__S (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__S (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__S (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__B2 (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A3 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__A3 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A3 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A3 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__A3 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__A3 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__A3 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09020__A (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__A (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__A (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__A2 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__A2 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__A2 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__B (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__S (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__S (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__A (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__A2 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__A2 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__A2 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__A2 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__A2 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__A2 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__A2 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__A2 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__S (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__S (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__S (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__S (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__S (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__S (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__A0 (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__A0 (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__A0 (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A0 (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A0 (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__A0 (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__A0 (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07732__A0 (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07677__A0 (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__A0 (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__A (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09480__A (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08830__A (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__A (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08491__A (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__A (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__A (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__A (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__A (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__A (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07677__S (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__S (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__S (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__S (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__A1 (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__A1 (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__A1 (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__A1 (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__A1 (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08022__A1 (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__A1 (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__A1 (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__A1 (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07695__A1 (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__S (.DIODE(_02598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__S (.DIODE(_02598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__S (.DIODE(_02598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07695__S (.DIODE(_02598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A1 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__A1 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A1 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__A1 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A1 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__A1 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A1 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__A1 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__A1 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__A1 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08383__A1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__A1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__A1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__A1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__A1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__A1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__A1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__A1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__A1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__A1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__A1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__A1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__A1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__A1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__S (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__S (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__S (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__S (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08416__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__A (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__A (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__A (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__A (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__A (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__B1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__B1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08420__B1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__B1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__B1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__B1 (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__B1 (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__B1 (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__B (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__A0 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__A0 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__A0 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__A0 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__A0 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A0 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A0 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A0 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__A0 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A0 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__S (.DIODE(_02648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__S (.DIODE(_02648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__S (.DIODE(_02648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__S (.DIODE(_02648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__A0 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__A0 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__A0 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A0 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__A0 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A0 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A0 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A0 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__A0 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__A0 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A0 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__A0 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__A0 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A0 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__A0 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A0 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__A0 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A0 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A0 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A0 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__S (.DIODE(_02659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__S (.DIODE(_02659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__S (.DIODE(_02659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__S (.DIODE(_02659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__B1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__B1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__B1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08840__B1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__B1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__B1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__B1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__B1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__B1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__S (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__S (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__S (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__S (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07854__S (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__S (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__S (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__S (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__B1 (.DIODE(_02714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__B1 (.DIODE(_02714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__B1 (.DIODE(_02714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__B1 (.DIODE(_02714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__B1 (.DIODE(_02714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__B1 (.DIODE(_02714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__B1 (.DIODE(_02714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__B1 (.DIODE(_02714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__B1 (.DIODE(_02714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__B1 (.DIODE(_02714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__S (.DIODE(_02717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__S (.DIODE(_02717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__S (.DIODE(_02717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__S (.DIODE(_02717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__B1 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__B1 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__B1 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__B1 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__B1 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__B1 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__B1 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__B1 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__B1 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07907__B1 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A2 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__A2 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A2 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__B1 (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__S (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__S (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__S (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__S (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__S (.DIODE(_02775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__S (.DIODE(_02775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__S (.DIODE(_02775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__S (.DIODE(_02775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__A0 (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08245__A0 (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__A0 (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A0 (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__A0 (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A0 (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__A0 (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__A0 (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__A0 (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__A0 (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__S (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__S (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__S (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08022__S (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A1 (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__A1 (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__A1 (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__A1 (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A1 (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__A1 (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__A1 (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08159__A1 (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A1 (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A1 (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__B1 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__B1 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__B1 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__B1 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__B1 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08722__B1 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__B1 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__B1 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__B1 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__B1 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__A1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__C1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09193__C1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08922__C1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__C1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__C1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__C1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__C1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__C1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__C1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__C1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A2 (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A2 (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__A2 (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__B (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__C1 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__C1 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__C1 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__C1 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__C1 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__C1 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__C1 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__C1 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__C1 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__C1 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__A0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__A0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__A0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08239__A0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__A0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__A0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__A0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__A0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A0 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__A0 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__A0 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__A0 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__A0 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__A0 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A0 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__A0 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__A0 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__A0 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A0 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A0 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__A0 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__A0 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__A0 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__A0 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A0 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A0 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A0 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__A0 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08545__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08418__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08712__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08546__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08199__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__S (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__S (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__S (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__S (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08418__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__A2 (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__A2 (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A2 (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__B1 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__B1 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__B1 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08804__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08789__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08622__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__A0 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__A0 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08563__A0 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__A0 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__A0 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08459__A0 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__A0 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A0 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__A0 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__A0 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__B1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__B1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__B1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__B1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__B1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08686__B1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__B1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__B1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__B1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__B1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__S (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__S (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__S (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__S (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08686__A1 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__A1 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A1 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A1 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A1 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__A1 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__A1 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__A1 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08416__A1 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__A1 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__A (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__A0 (.DIODE(_03103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__A0 (.DIODE(_03103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__A0 (.DIODE(_03109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__A0 (.DIODE(_03109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__A0 (.DIODE(_03109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A0 (.DIODE(_03109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08623__A0 (.DIODE(_03109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__A0 (.DIODE(_03109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__A0 (.DIODE(_03109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08502__A0 (.DIODE(_03109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A0 (.DIODE(_03109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__A0 (.DIODE(_03109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__A0 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__A0 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__A0 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08637__A0 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__A0 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__A0 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__A0 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08504__A0 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__A0 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__A0 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A0 (.DIODE(_03118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08727__A0 (.DIODE(_03118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A0 (.DIODE(_03118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08639__A0 (.DIODE(_03118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08627__A0 (.DIODE(_03118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__A0 (.DIODE(_03118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__A0 (.DIODE(_03118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__A0 (.DIODE(_03118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__A0 (.DIODE(_03118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__A0 (.DIODE(_03118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__A1 (.DIODE(_03141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__A1 (.DIODE(_03141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__A1 (.DIODE(_03141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08545__A1 (.DIODE(_03141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__A1 (.DIODE(_03141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__A1 (.DIODE(_03141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__A1 (.DIODE(_03141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__A1 (.DIODE(_03141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A1 (.DIODE(_03141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__A1 (.DIODE(_03141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__A (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09589__A (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__A (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__A (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__A (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__A (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08862__A (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08693__A (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__A (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A1 (.DIODE(_03169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__A1 (.DIODE(_03169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__A1 (.DIODE(_03169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A1 (.DIODE(_03169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__A1 (.DIODE(_03169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08864__A1 (.DIODE(_03169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08713__A1 (.DIODE(_03169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__A1 (.DIODE(_03169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__A1 (.DIODE(_03169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__A1 (.DIODE(_03169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__S (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__S (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__S (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__S (.DIODE(_03170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__A1 (.DIODE(_03172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__A1 (.DIODE(_03172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__A1 (.DIODE(_03172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__A1 (.DIODE(_03172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A1 (.DIODE(_03172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__A1 (.DIODE(_03172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__A1 (.DIODE(_03172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__A1 (.DIODE(_03172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08549__A1 (.DIODE(_03172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A1 (.DIODE(_03172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08887__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__S (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__S (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08549__S (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__S (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__A2 (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__A2 (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__A2 (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__B (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__A0 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09113__A0 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__A0 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__A0 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__A0 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__A0 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__A0 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__A0 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__A0 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__A0 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__A0 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08920__A1 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__A1 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08914__A1 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__A1 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__A1 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08853__A1 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__A1 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__A1 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__A1 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08690__A1 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__S (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__S (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__S (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__S (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__S (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__S (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__S (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08713__S (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__B1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__B1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__B1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__B1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__B1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__B1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08914__B1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08853__B1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__B1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__B1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__B1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__B1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__B1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__B1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__B1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__B1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__B1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__B1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__B1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__A2 (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A2 (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A2 (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__B (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08774__A (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A0 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A0 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09155__A0 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__A0 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__A0 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__A0 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08893__A0 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A0 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__A0 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__A0 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__A0 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A0 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09157__A0 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A0 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__A0 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__A0 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__A0 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__A0 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__A0 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__A0 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A0 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__A0 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__A0 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A0 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__A0 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A0 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__A0 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A0 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__A0 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__A0 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__S (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__S (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__S (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__S (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__B1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__B1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__B1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__B1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__B1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__B1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__B1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__B1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__B1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__B1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__S (.DIODE(_03388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__S (.DIODE(_03388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__S (.DIODE(_03388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__S (.DIODE(_03388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__A2 (.DIODE(_03440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A2 (.DIODE(_03440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A2 (.DIODE(_03440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__B (.DIODE(_03440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08940__A (.DIODE(_03451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__A (.DIODE(_03455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08950__A (.DIODE(_03459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A0 (.DIODE(_03461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A0 (.DIODE(_03461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__A0 (.DIODE(_03461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__A0 (.DIODE(_03461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A0 (.DIODE(_03461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A0 (.DIODE(_03461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A0 (.DIODE(_03461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__A0 (.DIODE(_03461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__A0 (.DIODE(_03461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__A0 (.DIODE(_03461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A1 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A1 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__A1 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__A1 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A1 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A1 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A1 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__A1 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__A1 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__A1 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A2 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A2 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__A2 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__A2 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A2 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A2 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A2 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__A2 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__A2 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__A2 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A3 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A3 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__A3 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__A3 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A3 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A3 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A3 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__A3 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__A3 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__A3 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__A0 (.DIODE(_03466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A0 (.DIODE(_03466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A0 (.DIODE(_03466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__A0 (.DIODE(_03466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A0 (.DIODE(_03466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A0 (.DIODE(_03466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__A0 (.DIODE(_03466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A0 (.DIODE(_03466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__A0 (.DIODE(_03466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A0 (.DIODE(_03466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__A1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__A1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__A1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__A1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__A2 (.DIODE(_03468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A2 (.DIODE(_03468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A2 (.DIODE(_03468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__A2 (.DIODE(_03468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A2 (.DIODE(_03468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A2 (.DIODE(_03468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__A2 (.DIODE(_03468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A2 (.DIODE(_03468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__A2 (.DIODE(_03468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A2 (.DIODE(_03468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__A3 (.DIODE(_03469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A3 (.DIODE(_03469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A3 (.DIODE(_03469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__A3 (.DIODE(_03469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A3 (.DIODE(_03469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A3 (.DIODE(_03469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__A3 (.DIODE(_03469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A3 (.DIODE(_03469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__A3 (.DIODE(_03469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A3 (.DIODE(_03469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__A2 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A2 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__A2 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A2 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__A2 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A2 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A2 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A2 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__A2 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__A2 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__A3 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A3 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__A3 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A3 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__A3 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A3 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A3 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A3 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__A3 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__A3 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__A0 (.DIODE(_03478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__A0 (.DIODE(_03478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__A0 (.DIODE(_03478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A0 (.DIODE(_03478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A0 (.DIODE(_03478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A0 (.DIODE(_03478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__A0 (.DIODE(_03478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__A0 (.DIODE(_03478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__A0 (.DIODE(_03478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__A0 (.DIODE(_03478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__A1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__A1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__A1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__A1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__A1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__A1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__A1 (.DIODE(_03479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__A2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__A2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__A2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__A2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__A2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__A2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__A2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__A3 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__A3 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__A3 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A3 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A3 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A3 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__A3 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__A3 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__A3 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__A3 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__A0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__A0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__A0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09029__A (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__A0 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A0 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__A0 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__A0 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A0 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__A0 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A0 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A0 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__A0 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08984__A0 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09030__A (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__A (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__A1 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A1 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__A1 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__A1 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A1 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__A1 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A1 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A1 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__A1 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08984__A1 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A2 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A2 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__A2 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A2 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A2 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__A2 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__A2 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A2 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09031__A (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__A (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__A2 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A2 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__A2 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__A2 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A2 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__A2 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A2 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A2 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__A2 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08984__A2 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A3 (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A3 (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__A3 (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A3 (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A3 (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__A3 (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__A3 (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A3 (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09032__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__A3 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A3 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__A3 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__A3 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A3 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__A3 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A3 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A3 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__A3 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08984__A3 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A0 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A0 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__A0 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A0 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A0 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__A0 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__A0 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A0 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A0 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__A (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__A0 (.DIODE(_03494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A0 (.DIODE(_03494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__A0 (.DIODE(_03494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__A0 (.DIODE(_03494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__A0 (.DIODE(_03494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A0 (.DIODE(_03494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A0 (.DIODE(_03494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A0 (.DIODE(_03494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09060__A0 (.DIODE(_03494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A0 (.DIODE(_03494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A1 (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A1 (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__A1 (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A1 (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A1 (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__A1 (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__A1 (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A1 (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A1 (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__A (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__A1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__A1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__A1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__A1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09060__A1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A2 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A2 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__A2 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A2 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A2 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__A2 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__A2 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A2 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A2 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__A (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09060__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A3 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A3 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__A3 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A3 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A3 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__A3 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__A3 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A3 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A3 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__A (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__A3 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A3 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__A3 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__A3 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__A3 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A3 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A3 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A3 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09060__A3 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A3 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__A0 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A0 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A0 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__A0 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A0 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A0 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A0 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A0 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__A0 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A0 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__A1 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A1 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A1 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__A1 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A1 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A1 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A1 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A1 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__A1 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A1 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__A2 (.DIODE(_03505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A2 (.DIODE(_03505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A2 (.DIODE(_03505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__A2 (.DIODE(_03505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A2 (.DIODE(_03505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A2 (.DIODE(_03505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A2 (.DIODE(_03505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A2 (.DIODE(_03505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__A2 (.DIODE(_03505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A2 (.DIODE(_03505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__A3 (.DIODE(_03506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A3 (.DIODE(_03506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A3 (.DIODE(_03506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__A3 (.DIODE(_03506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A3 (.DIODE(_03506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A3 (.DIODE(_03506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A3 (.DIODE(_03506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A3 (.DIODE(_03506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__A3 (.DIODE(_03506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A3 (.DIODE(_03506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A0 (.DIODE(_03511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__A0 (.DIODE(_03511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A0 (.DIODE(_03511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__A0 (.DIODE(_03511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__A0 (.DIODE(_03511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A0 (.DIODE(_03511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A0 (.DIODE(_03511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A0 (.DIODE(_03511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__A0 (.DIODE(_03511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__A0 (.DIODE(_03511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A1 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__A1 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A1 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__A1 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__A1 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A1 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A1 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A1 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__A1 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__A1 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A2 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__A2 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A2 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__A2 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__A2 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A2 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A2 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A2 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__A2 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__A2 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A3 (.DIODE(_03514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__A3 (.DIODE(_03514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A3 (.DIODE(_03514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__A3 (.DIODE(_03514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__A3 (.DIODE(_03514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A3 (.DIODE(_03514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A3 (.DIODE(_03514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A3 (.DIODE(_03514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__A3 (.DIODE(_03514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__A3 (.DIODE(_03514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A0 (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A0 (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09724__A0 (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__A0 (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__A0 (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A0 (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__A0 (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A0 (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A0 (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__A0 (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09724__A1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__A1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__A1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__A1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__A1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09724__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A3 (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A3 (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09724__A3 (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__A3 (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__A3 (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A3 (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__A3 (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A3 (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A3 (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__A3 (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__A1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__A1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__A1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__A1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A2 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__A2 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A2 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A2 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A2 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__A2 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__A2 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A2 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A2 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__A2 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A3 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__A3 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A3 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A3 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A3 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__A3 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__A3 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A3 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A3 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__A3 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A2 (.DIODE(_03530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__A0 (.DIODE(_03530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__A0 (.DIODE(_03530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__A0 (.DIODE(_03530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A0 (.DIODE(_03530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A0 (.DIODE(_03530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A0 (.DIODE(_03530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A0 (.DIODE(_03530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__A0 (.DIODE(_03530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__A0 (.DIODE(_03530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__B (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__B (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__B (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__B (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__A0 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__A2 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A2 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A2 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__A2 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__A2 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A2 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__A2 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A2 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A2 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__A1 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__A3 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A3 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A3 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__A3 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__A3 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__A0 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A0 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__A0 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A0 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A0 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__A0 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__A0 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A0 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__A0 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A0 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__A1 (.DIODE(_03537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A1 (.DIODE(_03537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__A1 (.DIODE(_03537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A1 (.DIODE(_03537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A1 (.DIODE(_03537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__A1 (.DIODE(_03537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__A1 (.DIODE(_03537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A1 (.DIODE(_03537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__A1 (.DIODE(_03537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A1 (.DIODE(_03537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__A2 (.DIODE(_03538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A2 (.DIODE(_03538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__A2 (.DIODE(_03538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A2 (.DIODE(_03538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A2 (.DIODE(_03538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__A2 (.DIODE(_03538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__A2 (.DIODE(_03538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A2 (.DIODE(_03538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__A2 (.DIODE(_03538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A2 (.DIODE(_03538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__A3 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A3 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__A3 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A3 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A3 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__A3 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__A3 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A3 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__A3 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A3 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__A0 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A0 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__A0 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__A0 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A0 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A0 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__A0 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__A0 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__A0 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__A0 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__A1 (.DIODE(_03542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A1 (.DIODE(_03542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__A1 (.DIODE(_03542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__A1 (.DIODE(_03542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A1 (.DIODE(_03542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A1 (.DIODE(_03542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__A1 (.DIODE(_03542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__A1 (.DIODE(_03542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__A1 (.DIODE(_03542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__A1 (.DIODE(_03542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__A3 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A3 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__A3 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__A3 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A3 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A3 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__A3 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__A3 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__A3 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__A3 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A0 (.DIODE(_03546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09886__A0 (.DIODE(_03546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__A0 (.DIODE(_03546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A0 (.DIODE(_03546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__A0 (.DIODE(_03546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__A0 (.DIODE(_03546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__A0 (.DIODE(_03546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A0 (.DIODE(_03546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A0 (.DIODE(_03546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A0 (.DIODE(_03546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09886__A1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__A1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__A1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__A1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__A1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09886__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A3 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09886__A3 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__A3 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A3 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__A3 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__A3 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__A3 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A3 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A3 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A3 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09113__S (.DIODE(_03592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__S (.DIODE(_03592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__S (.DIODE(_03592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__S (.DIODE(_03592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__S (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__A0 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__A0 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A0 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__A0 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A0 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__A0 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A0 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__A0 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__A0 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__A0 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__S (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__S (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09157__S (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09155__S (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__A1 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__A1 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__A1 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__A1 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A1 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A1 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__A1 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09191__A1 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__A1 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__A1 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__S (.DIODE(_03677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__S (.DIODE(_03677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__S (.DIODE(_03677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__S (.DIODE(_03677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__A0 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__A2 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__A0 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__A0 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A0 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__A0 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__A0 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__A0 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A0 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A0 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__A1 (.DIODE(_03698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__A1 (.DIODE(_03698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A1 (.DIODE(_03698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__A1 (.DIODE(_03698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A1 (.DIODE(_03698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__A1 (.DIODE(_03698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__A1 (.DIODE(_03698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__A1 (.DIODE(_03698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A1 (.DIODE(_03698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A1 (.DIODE(_03698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__A2 (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__A2 (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__A2 (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__B1 (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__B1 (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__B1 (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A0 (.DIODE(_03749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A0 (.DIODE(_03749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__A2 (.DIODE(_03758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__A2 (.DIODE(_03758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__A2 (.DIODE(_03758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A0 (.DIODE(_03758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A2 (.DIODE(_03758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A1 (.DIODE(_03758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A0 (.DIODE(_03758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A2 (.DIODE(_03758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__A2 (.DIODE(_03758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A0 (.DIODE(_03758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__A3 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__A3 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__A3 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A1 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A3 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A0 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A1 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A3 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__A3 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A1 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__A0 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__A0 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__A0 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A2 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A0 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A3 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A2 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A0 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__A0 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A2 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__A1 (.DIODE(_03761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__A1 (.DIODE(_03761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__A1 (.DIODE(_03761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A3 (.DIODE(_03761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A1 (.DIODE(_03761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A2 (.DIODE(_03761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A3 (.DIODE(_03761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A1 (.DIODE(_03761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__A1 (.DIODE(_03761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A3 (.DIODE(_03761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A0 (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A0 (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A0 (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A0 (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__A0 (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__A0 (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__A0 (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__A0 (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__A0 (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A0 (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A2 (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A2 (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A2 (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A2 (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__A2 (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__A2 (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__A2 (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__A2 (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__A2 (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A2 (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A3 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A3 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A3 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A3 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__A3 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__A3 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__A3 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__A3 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__A3 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A3 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__B (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10173__A0 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A0 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__A2 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__A2 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__A2 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A2 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__A2 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__A2 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A2 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__A2 (.DIODE(_03787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10173__A1 (.DIODE(_03787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A1 (.DIODE(_03787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__A3 (.DIODE(_03787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__A3 (.DIODE(_03787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__A3 (.DIODE(_03787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A3 (.DIODE(_03787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__A3 (.DIODE(_03787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__A3 (.DIODE(_03787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A3 (.DIODE(_03787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__A0 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A0 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__A0 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__A0 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__A0 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__A0 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A0 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A0 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__A0 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A0 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__A1 (.DIODE(_03807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A1 (.DIODE(_03807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__A1 (.DIODE(_03807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__A1 (.DIODE(_03807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__A1 (.DIODE(_03807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__A1 (.DIODE(_03807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A1 (.DIODE(_03807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A1 (.DIODE(_03807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__A1 (.DIODE(_03807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A1 (.DIODE(_03807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__A2 (.DIODE(_03808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A2 (.DIODE(_03808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__A2 (.DIODE(_03808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__A2 (.DIODE(_03808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__A2 (.DIODE(_03808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__A2 (.DIODE(_03808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A2 (.DIODE(_03808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A2 (.DIODE(_03808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__A2 (.DIODE(_03808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A2 (.DIODE(_03808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__A3 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A3 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__A3 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__A3 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__A3 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__A3 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A3 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A3 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__A3 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A3 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__A0 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A0 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A0 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__A0 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A0 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__A0 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__A0 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__A0 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__A0 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A0 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A1 (.DIODE(_03817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__A2 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A2 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A2 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__A2 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A2 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__A2 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__A2 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__A2 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__A2 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A2 (.DIODE(_03818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__A3 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A3 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A3 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__A3 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A3 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__A3 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__A3 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__A3 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__A3 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A3 (.DIODE(_03819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A0 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__A0 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__A0 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__A0 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09718__A0 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__A0 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A0 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A0 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__A0 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__A0 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__S (.DIODE(_03870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A0 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__A0 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__A0 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A0 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__A0 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__A0 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__A0 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__A0 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__A0 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A0 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__A0 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09837__A0 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__A0 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__A0 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__A0 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__A0 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__A0 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__A0 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__A0 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__A0 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__S (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__S (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__S (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__S (.DIODE(_03881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__A1 (.DIODE(_03914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__S (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__S (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__S (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__S (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09556__S (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__S (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__S (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__S (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__S (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__S (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__S (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__S (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__A1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10069__A1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__A1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__A1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__A1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__A1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__A1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09796__A1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__A1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__A1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A2 (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A2 (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__A2 (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__B (.DIODE(_03990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__C (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__C (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__C (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__C (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__C (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__C (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__C (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__C (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__S (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__S (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09686__A2 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__S (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__S (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__S (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09718__S (.DIODE(_04106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__S (.DIODE(_04130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__S (.DIODE(_04130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__S (.DIODE(_04130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__S (.DIODE(_04130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__S (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__S (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__S (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__S (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__S (.DIODE(_04171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__S (.DIODE(_04171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__S (.DIODE(_04171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__S (.DIODE(_04171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10125__A1 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__A1 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__A1 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__A1 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__A1 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__A1 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10047__A1 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A1 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10039__A1 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__A1 (.DIODE(_04181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09830__S (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__S (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__S (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__S (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A0 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A0 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A0 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A0 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__A0 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__A0 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__A0 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__A0 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__A0 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A0 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A1 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A1 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A1 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A1 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__A1 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__A1 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__A1 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__A1 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__A1 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A1 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A2 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A2 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A2 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A2 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__A2 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__A2 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__A2 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__A2 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__A2 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A2 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A3 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A3 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A3 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A3 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__A3 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__A3 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__A3 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__A3 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__A3 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A3 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__S (.DIODE(_04340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__S (.DIODE(_04340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__S (.DIODE(_04340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__S (.DIODE(_04340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10020__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__S (.DIODE(_04374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__S (.DIODE(_04374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__S (.DIODE(_04374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__S (.DIODE(_04374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__S (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__S (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__S (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__S (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__S (.DIODE(_04398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__S (.DIODE(_04398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__S (.DIODE(_04398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__S (.DIODE(_04398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10388__A (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__A (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__A (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__A (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__A (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__A (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__A (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__A1 (.DIODE(_04417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__A (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10393__A (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__A (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10350__A (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__A (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10309__A (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__A (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10266__A (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__A (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10132__A1 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A2 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__A2 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__A2 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__B (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__B1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__B1 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__B1 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__B1 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__B1 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__A (.DIODE(_04554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A (.DIODE(_04554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__A (.DIODE(_04554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__A (.DIODE(_04554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__A (.DIODE(_04554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__A (.DIODE(_04554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__A (.DIODE(_04554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A (.DIODE(_04554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A (.DIODE(_04554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__A (.DIODE(_04554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10430__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10389__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10396__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__A (.DIODE(_04622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A (.DIODE(_04622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__A (.DIODE(_04622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__A (.DIODE(_04622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__A (.DIODE(_04622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__A (.DIODE(_04622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10429__A (.DIODE(_04622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__A (.DIODE(_04622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__A (.DIODE(_04622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__A (.DIODE(_04622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10524__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10535__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10454__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__A (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__A (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10574__A (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__A (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10539__A (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10531__A (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__A (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__A (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__A (.DIODE(_04738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A (.DIODE(_04738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A (.DIODE(_04738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__A (.DIODE(_04738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10620__A (.DIODE(_04738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__A (.DIODE(_04738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__A (.DIODE(_04738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__A (.DIODE(_04738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__A (.DIODE(_04738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__A (.DIODE(_04738_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2930_A (.DIODE(\c.cfg_i_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06975__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04855__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04850__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04814__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06311__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04969__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04863__B (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04860__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04829__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06319__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05286__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04927__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04877__B (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04875__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04838__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__C (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09465__C (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__C (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__C (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__C (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__C (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06271__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05150__C (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04995__A (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04817__B (.DIODE(\c.genblk1.genblk1.subs.c0.cfg_i_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__B1 (.DIODE(\c.genblk1.genblk1.subs.c0.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__A_N (.DIODE(\c.genblk1.genblk1.subs.c0.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__A_N (.DIODE(\c.genblk1.genblk1.subs.c0.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__C (.DIODE(\c.genblk1.genblk1.subs.c0.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__C (.DIODE(\c.genblk1.genblk1.subs.c0.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08762__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06076__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05992__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05907__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08762__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06079__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05992__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05623__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06079__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05907__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05626__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05901__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05631__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05903__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05631__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08762__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05992__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05907__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05629__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05630__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__C1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06571__C1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06244__C1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06072__C1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05897__C1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05712__C1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05618__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.grst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14351__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14355__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14359__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06021__S (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06016__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06015__C1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4096_A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06008__S (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06005__S (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06003__S0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06001__S0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06000__S0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.lut_in_sels[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04907__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.rst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04855__B (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.rst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04842__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.rst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04824__A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.luts.rst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14346__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14567__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14571__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14575__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.imuxs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14562__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold523_A (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05869__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05857__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05839__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05827__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14783__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14778__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A0 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14995__D (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__A3 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A2 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A1 (.DIODE(\c.genblk1.genblk1.subs.c0.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__B1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__A_N (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__A_N (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__C (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__C (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10523__B1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__B (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__B (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__A_N (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__A_N (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__A (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__A (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07371__A (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__A (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__A (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__A (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__D (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13472__D (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__B1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__B (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__B (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__A_N (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__A_N (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13688__D (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13904__D (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14121__D (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[1].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__B1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__A_N (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__A_N (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06298__C (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06272__C (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06481__A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06579__A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06482__A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3044_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06449__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06430__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06423__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06403__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3099_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06454__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06434__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06418__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06411__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3039_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06459__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06431__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06424__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06404__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3074_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06445__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06433__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06421__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06406__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__D (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2959_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06550__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06538__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06525__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06512__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2961_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06545__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06533__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06521__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06499__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2978_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06539__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06526__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06504__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2960_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06544__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06536__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06517__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06509__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3308_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1927_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__D (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06578__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3083_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06638__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06610__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06590__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3045_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06643__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06622__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06606__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06596__A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__D (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06674__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3079_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06732__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06711__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06698__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3029_A (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06685__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.ibufs[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13255__D (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06763__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[2].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__B1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__A_N (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__A_N (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04817__C (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05814__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06265__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06262__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06162__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05721__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05725__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05726__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05816__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05720__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05817__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05722__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05727__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A3 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05728__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.globs[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2947_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05693__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05673__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05658__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05639__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3100_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05679__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05670__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05652__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05641__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__D (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.imuxs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2025_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2832_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.luts.ram[2][30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__D (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__B (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[0].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3067_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05784__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05768__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05761__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05748__B (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3108_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05785__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05770__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05763__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05739__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3070_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05787__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05772__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05755__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05743__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4035_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05752__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05750__A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05741__C1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05736__C1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.lut_in_sels[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2842_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[0][31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1891_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2083_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1608_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold639_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[1][31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2886_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2115_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1680_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1032_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.luts.ram[2][31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11956__D (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__A1 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10172__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05815__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[1].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2924_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06145__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06122__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06107__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06088__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2918_A (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06131__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06119__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06101__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06090__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.ibufs[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__D (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.imuxs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__D (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06261__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06161__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[2].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__D (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.imuxs[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__D (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06267__A2 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06247__A0 (.DIODE(\c.genblk1.genblk1.subs.cs[3].c.genblk1.genblk1.leaf.lbs[3].lb_.o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__B1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04996__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04817__A_N (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4142_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04896__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04912__A0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4112_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04937__A0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__B2 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04939__A0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09060__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04949__A0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4164_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09060__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4103_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09061__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09056__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4086_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4058_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4138_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04869__B2 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4121_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__A_N (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__B1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[0].x.selects.o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__B1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05150__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04996__A_N (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05045__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4082_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05070__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05086__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05103__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4122_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4098_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3806_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[37] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09320__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[37] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__A_N (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[37] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3972_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__A2 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__A2 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[38] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3942_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__C1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05025__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4095_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[1].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__B1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05305__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05150__A_N (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05201__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4081_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4060_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09628__A_N (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__C1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4066_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09628__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4167_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05179__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05183__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[2].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__B1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05463__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05305__A_N (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.cfgd ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4127_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05382__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4068_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__A_N (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__C1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4028_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4171_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4160_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05400__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05417__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3878_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__A_N (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__C1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4007_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4050_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4021_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__B1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3790_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4026_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09886__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4169_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09886__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__B (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09988__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05321__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05338__A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4071_A (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.dns[3].x.selects.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold161_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3071_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2940_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold183_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__S (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10193__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05494__A0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4055_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__B2 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__B1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3961_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__S (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__C1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3971_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__S (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4004_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4072_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__A1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4148_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__S (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3974_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__B1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10216__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__S1 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4076_A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__S0 (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__S (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10204__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__A (.DIODE(\c.genblk1.genblk1.subs.sw.up.x.selects.o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(cfg));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold15_A (.DIODE(cfg_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold7_A (.DIODE(cfg_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold6_A (.DIODE(cfg_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold18_A (.DIODE(cfg_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold8_A (.DIODE(cfg_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1_A (.DIODE(grst));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3_A (.DIODE(m[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold14_A (.DIODE(m[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold40_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(up_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(up_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(up_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(up_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(up_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(up_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(up_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(up_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(up_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(up_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(up_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(up_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(up_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(up_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(up_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(up_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__C (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__C (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__A0 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A0 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09367__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__08997__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__A3 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09040__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__A3 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__A3 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__A3 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09042__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09010__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09011__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09012__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__08980__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A3 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08982__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09035__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__05463__A_N (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__14340__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14343__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14207__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14214__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14167__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14262__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14168__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14301__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14254__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14215__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14317__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14270__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14223__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13957__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14366__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14176__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14160__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14357__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14354__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14356__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14351__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14355__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14363__CLK (.DIODE(clknet_leaf_18_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11105__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11099__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11137__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11097__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__CLK (.DIODE(clknet_leaf_56_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11516__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11522__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11070__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11109__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11107__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__CLK (.DIODE(clknet_leaf_59_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10844__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11085__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14346__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14778__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14562__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14995__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__CLK (.DIODE(clknet_leaf_63_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10989__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11084__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11124__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__CLK (.DIODE(clknet_leaf_64_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__15017__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10820__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10704__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10740__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10744__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10725__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10808__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10810__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__15016__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__15023__CLK (.DIODE(clknet_leaf_65_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14714__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14781__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14976__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14780__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14996__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14563__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14349__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14348__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14977__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14779__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14930__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14883__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14979__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14347__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10845__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10709__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10826__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10858__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10856__CLK (.DIODE(clknet_leaf_67_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11357__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11302__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__CLK (.DIODE(clknet_leaf_80_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12180__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12188__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12136__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__CLK (.DIODE(clknet_leaf_102_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12381__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12373__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12324__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12231__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12174__CLK (.DIODE(clknet_leaf_115_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12667__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__CLK (.DIODE(clknet_leaf_126_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12721__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12622__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12582__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12612__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__CLK (.DIODE(clknet_leaf_134_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12692__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12684__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12688__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12696__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__CLK (.DIODE(clknet_leaf_137_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13572__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13883__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13836__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13897__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13573__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13581__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13583__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13899__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13900__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13764__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13717__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13901__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13902__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13797__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13844__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13840__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13746__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13891__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13903__CLK (.DIODE(clknet_leaf_175_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14150__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13994__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14040__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13946__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14039__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14086__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13993__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14087__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14129__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14127__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14128__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14132__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13947__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14041__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14042__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14088__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13948__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14133__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14089__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13740__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13787__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13995__CLK (.DIODE(clknet_leaf_190_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_clk_A (.DIODE(clknet_1_0_1_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_clk_A (.DIODE(clknet_1_0_1_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_clk_A (.DIODE(clknet_1_1_1_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_clk_A (.DIODE(clknet_1_1_1_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_clk_A (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_clk_A (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_clk_A (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_clk_A (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_clk_A (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_clk_A (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_clk_A (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_clk_A (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_190_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_1_0_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_188_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_187_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_2_0_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_186_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_185_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_184_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_183_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_182_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_181_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_180_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_179_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_178_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_177_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_176_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_175_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_174_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_173_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_172_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_171_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_170_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_169_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_168_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_3_0_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_161_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_160_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_159_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_158_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_157_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_156_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_155_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_154_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_153_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_152_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_151_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_150_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_149_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_167_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_166_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_165_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_164_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_163_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_162_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_125_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_124_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_123_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_122_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_121_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_148_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_147_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_146_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_145_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_144_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_143_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_142_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_141_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_140_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_139_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_138_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_136_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_137_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_135_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_134_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_133_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_132_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_131_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_130_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_129_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_128_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_127_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_126_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_119_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__D (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__D (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__D (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__D (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__D (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__D (.DIODE(net1716));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__D (.DIODE(net1927));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__D (.DIODE(net1963));
 sky130_fd_sc_hd__diode_2 ANTENNA__11668__D (.DIODE(net2061));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__D (.DIODE(net2119));
 sky130_fd_sc_hd__diode_2 ANTENNA__11925__D (.DIODE(net2151));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__D (.DIODE(net2868));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__D (.DIODE(net2878));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__D (.DIODE(net2922));
 sky130_fd_sc_hd__diode_2 ANTENNA__14144__D (.DIODE(net2966));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__D (.DIODE(net3107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__A (.DIODE(net3415));
 sky130_fd_sc_hd__diode_2 ANTENNA__09279__B1 (.DIODE(net3415));
 sky130_fd_sc_hd__diode_2 ANTENNA__04854__B2 (.DIODE(net3415));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__A2 (.DIODE(net3826));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__A1 (.DIODE(net3826));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__A (.DIODE(net3826));
 sky130_fd_sc_hd__diode_2 ANTENNA__05440__A1 (.DIODE(net3826));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A (.DIODE(net3890));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__B1 (.DIODE(net3890));
 sky130_fd_sc_hd__diode_2 ANTENNA__05391__A (.DIODE(net3890));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__A0 (.DIODE(net4071));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1064 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1265 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1255 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1215 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1256 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1256 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1258 ();
 assign io_o = net36;
endmodule

